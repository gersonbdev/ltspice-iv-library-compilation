SCN14
.OPTIONS LIMPTS=1000
*SPICE_NET
*INCLUDE SCN.LIB
.AC DEC 10 1K 10MEG
*ALIAS  V(19)=VOUT
.PRINT AC  V(19)  VP(19) 
R73 2 3 100.86K
R74 19 5 25.42K
R75 6 5 17.72K
R76 7 5 11.52K
V14 3 0 AC 1
R77 8 9 99.83K
R78 10 9 68.15K
R79 11 9 10.18K
R80 8 5 13.84K
R82 12 9 16.61K
R84 13 14 20.93K
R85 15 14 45.2K
R86 12 14 25.52K
R87 14 16 25.72K
R88 2 17 99.73K
R89 2 16 23.6K
R90 2 18 16.75K
X8 2 0 18 0 16 17 14 13 0 15 12 9 11 8 10 8 5 7 6 19 1 LT6410D 
V13 1 0 10
.END