SCN2
*SPICE_NET
*INCLUDE SCN.LIB
.AC DEC 50 1K 500K
.OPTIONS PIVTOL=1E-20 LIMPTS=20000
*.TRAN .05U 50U
*ALIAS  V(1)=VOUT
*ALIAS  V(20)=VOUT
.PRINT AC  V(1)  VP(1)  V(20)  VP(20) 
.PRINT TRAN  V(1)  V(20) 
X19 31 30 19 34 ZINT  {TD=1U C=32P } 
X2 35 36 2 33 ZINT  {TD=1U C=32P } 
X4 1 35 CRES  {C=2P } 
X5 5 35 CRES  {C=2P } 
X8 2 29 NSTR  {TD=1U C=2P } 
X9 28 29 1 32 ZINT  {TD=1U C=32P } 
E1 3 0 15 4 20K
X11 3 35 NSTR  {TD=1U C=2P } 
X20 20 31 CRES  {C=2P } 
X21 16 31 CRES  {C=2P } 
X22 19 38 NSTR  {TD=1U C=2P } 
X23 37 38 20 40 ZINT  {TD=1U C=32P } 
X24 18 31 NSTR  {TD=1U C=2P } 
E2 18 0 15 17 20K
C2 5 2 
.END