SCN13
.OPTIONS LIMPTS=1000
*SPICE_NET
*INCLUDE SCN.LIB
.AC DEC 100 1K 100K
*ALIAS  V(16)=VOUT
.PRINT AC  V(16)  VP(16) 
R12 12 14 46.95K
R14 15 20 10.5K
R15 16 20 39.42K
R16 17 20 13.19K
V2 14 0 AC 1
R17 1 5 10K
R18 3 5 70.3K
R19 2 5 16.3K
R20 1 20 17.9K
R21 2 20 69.7K
R22 4 5 27.46K
R23 7 5 6.9K
R24 7 8 10K
R25 6 8 81.5K
R26 4 8 14.72K
R27 8 25 93.93K
R28 12 10 11.81K
R29 12 25 38.25K
R30 12 11 10K
X2 12 0 11 0 25 10 8 7 0 6 4 5 2 0 3 1 20 17 16 15 9 LT6450D 
V1 9 0 2
.END