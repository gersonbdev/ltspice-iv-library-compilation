SCN9
*SPICE_NET
*INCLUDE SCN.LIB
*INCLUDE NONLIN.LIB
.AC LIN 200 1.5K 2.5K
.OPTIONS ACCT PIVTOL=1E-20 LIMPTS=1000
*ALIAS  V(13)=VOUT
*ALIAS  V(1)=VL1
*ALIAS  V(6)=VL2
.PRINT AC  V(13)  VP(13)  V(1)  VP(1) 
.PRINT AC  V(6)  VP(6) 
.PRINT TRAN  V(13)  V(1)  V(6) 
R21 3 2 5K
R31 3 5 152K
R41 3 1 5.27K
RL1 1 7 10.74K
V1 4 0 PULSE 0 1 AC 1
RH1 2 7 13.2K
R22 7 9 5.26K
R32 7 10 151.8K
R42 7 6 5K
X2 15 0 13 11 12 UA741
V2 12 0 -15
V3 11 0 15
RH2 9 15 5K
RG 15 13 37.3K
RL2 6 15 6.11K
VCLK 14 0 .4
*SET TO .4 FOR 2KHz NATURAL FREQUENCY 
*SET TO 1 FOR 500KHZ, GAIN = 100
*SET TO 4 FOR 20KHz NATURAL FREQUENCY 
C1 3 1 12P
C2 7 6 20P
X3 3 0 2 0 5 1 7 10 6 14 14 9 0 LT60L100 
R11 4 3 155.93K
.END