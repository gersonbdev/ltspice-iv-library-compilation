SCN7
*SPICE_NET
*INCLUDE SCN.LIB
.AC DEC 50 1K 500K
.OPTIONS ACCT LIMPTS=10000 PIVTOL=1E-20
.TRAN 20U 4M
*ALIAS  V(7)=VOUTA
*ALIAS  V(8)=VOUTB
.PRINT AC  V(7)  VP(7)  V(8)  VP(8) 
.PRINT TRAN  V(7)  V(8) 
R2 1 2 100K
R3 4 6 10K
R4 4 5 100K
V1 9 0 PULSE 0 2 AC 1
V2 10 0 1
V3 11 0 PULSE 0 2 AC 1
X3 1 0 3 11 2 7 4 5 8 10 10 6 9 MF10H100 
R1 1 3 10K
.END