IBIS
*SPICE_NET
.TRAN .1N 150N
*INCLUDE IBIS1.LIB
.SUBCKT PCIOB 100   4      300 400 500
*Connections    Input Output VCC VEE Enable
*Passed Parameters; Min
*dEFINE {RTF}=20K
*dEFINE {RTR}=20K
* Input Control
B1 820 0 V=V(100) & V(500)
B2 830 0 V= V(500) & ~V(100)
* Up and Down Ramps
B3 300 850 I= V(830) > 1.2   ? 0 : V(300,850) / 20K
B4 840 400 I= V(820) > 1.2 ? 0 : V(840,400) / 20K
C1 300 850 .01P
C2 840 400 .01P
S1 220 850 0 820 SMOD
S2 840 220 0 830 SMOD
.MODEL SMOD SW RON=.1M ROFF=1E15 VT=-1.2 VH=.1
G1 8 400 2 8 1
R1 6 400 1
G2 300 8 8 3 1
R2 300 6 1
* Pull-up/Pull-down structures; Max
XEPL_DN 2 400 8 840 EPWL_DNX
XEPL_UP 3 300 850 8 EPWL_UPX
* Diode Clamps
XVCC_OUT 6 300 300 6 VCC_OUT
XGND_OUT 6 400 6 400 GND_OUT
* Package Parasitics; Min
ROSNB 5 1 100
ROPKG 1 4 .100
COPKG 4 400 1.00P
CCOMP 5 400 4.00P
LOPKG 5 1 8.00N
* Voltage Sources for measuring currents
V5 6 5 
V6 8 6 
V7 220 8 
.ENDS
*Subcircuits for the IBIS1 Topology
.SUBCKT GND_OUT  3    4    1   2
*                OUT+ OUT- IN+ IN-
B1 3 4 I= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + -292.99998M :
+ (V(1,2) < -1.0000000) ? 66.999997M*V(1,2) + 41.999998M :
+ (V(1,2) < -899.99996M) ? 119.99999M*V(1,2) + 94.999995M :
+ (V(1,2) < -799.99996M) ? 69.999997M*V(1,2) + 49.999998M :
+ (V(1,2) < -699.99997M) ? 35.999998M*V(1,2) + 22.799999M :
+ (V(1,2) < -599.99997M) ? 11.999999M*V(1,2) + 5.9999997M :
+ (V(1,2) < -499.99998M) ? 6.9999997M*V(1,2) + 2.9999999M :
+ (V(1,2) < -399.99998M) ? 3.9999998M*V(1,2) + 1.4999999M :
+ (V(1,2) < 0.0000000E+00) ? 250.00000U*V(1,2) + -6.6174449E-12 :
+ 1.0000000N*V(1,2) + 0.0000000E+00
.ENDS
*
.SUBCKT VCC_OUT 3    4    1   2
*               OUT+ OUT- IN+ IN-
B1 3 4 I= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + 292.99999M :
+ (V(1,2) < -1.0000000) ? -66.999997M*V(1,2) + -41.999998M :
+ (V(1,2) < -899.99996M) ? -119.99999M*V(1,2) + -94.999995M :
+ (V(1,2) < -799.99996M) ? -69.999997M*V(1,2) + -49.999998M :
+ (V(1,2) < -699.99997M) ? -35.999998M*V(1,2) + -22.799999M :
+ (V(1,2) < -599.99997M) ? -11.999999M*V(1,2) + -5.9999997M :
+ (V(1,2) < -499.99998M) ? -6.9999997M*V(1,2) + -2.9999999M :
+ (V(1,2) < -399.99998M) ? -3.9999998M*V(1,2) + -1.4999999M :
+ (V(1,2) < 0.0000000E+00) ? -250.00000U*V(1,2) + 6.6174449E-12 :
+ 1.0000000N*V(1,2) + 0.0000000E+00
.ENDS
*
.SUBCKT EPWL_UPX 3    4    1   2
*                OUT+ OUT- IN+ IN-
B1 3 4 V= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + 137.00000M :
+ (V(1,2) < -4.0000000) ? -8.9999996M*V(1,2) + 91.999996M :
+ (V(1,2) < -3.0000000) ? -9.9999995M*V(1,2) + 87.999996M :
+ (V(1,2) < -2.0000000) ? -21.999999M*V(1,2) + 51.999998M :
+ (V(1,2) < -1.0000000) ? -31.999998M*V(1,2) + 31.999998M :
+ (V(1,2) < 0.0000000E+00) ? -63.999997M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 499.99998M) ? -75.999996M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 1.0000000) ? -51.999998M*V(1,2) + -11.999999M :
+ (V(1,2) < 1.5000000) ? -37.999998M*V(1,2) + -25.999999M :
+ (V(1,2) < 2.0000000) ? -25.999999M*V(1,2) + -43.999998M :
+ (V(1,2) < 2.5000000) ? -27.999999M*V(1,2) + -39.999998M :
+ (V(1,2) < 3.0000000) ? -15.999999M*V(1,2) + -69.999997M :
+ (V(1,2) < 3.5000000) ? -9.9999995M*V(1,2) + -87.999996M :
+ (V(1,2) < 4.0000000) ? -9.9999995M*V(1,2) + -87.999996M :
+ (V(1,2) < 4.5000000) ? -9.9999995M*V(1,2) + -87.999996M :
+ (V(1,2) < 5.0000000) ? -7.9999996M*V(1,2) + -96.999995M :
+ (V(1,2) < 10.0000000) ? -1.0000000M*V(1,2) + -131.99999M :
+ 1.0000000N*V(1,2) + -142.00000M
.ENDS
*
.SUBCKT EPWL_DNX  3    4    1   2
*                 OUT+ OUT- IN+ IN-
B1 3 4 V= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + -214.99998M :
+ (V(1,2) < -4.0000000) ? 2.9999999M*V(1,2) + -199.99999M :
+ (V(1,2) < -3.0000000) ? 4.9999998M*V(1,2) + -191.99999M :
+ (V(1,2) < -2.0000000) ? 18.999999M*V(1,2) + -149.99999M :
+ (V(1,2) < -1.0000000) ? 117.99999M*V(1,2) + 47.999998M :
+ (V(1,2) < 0.0000000E+00) ? 69.999997M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 499.99998M) ? 139.99999M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 1.0000000) ? 113.99999M*V(1,2) + 12.999999M :
+ (V(1,2) < 1.5000000) ? 73.999996M*V(1,2) + 52.999997M :
+ (V(1,2) < 2.0000000) ? 47.999998M*V(1,2) + 91.999996M :
+ (V(1,2) < 2.5000000) ? 29.999999M*V(1,2) + 127.99999M :
+ (V(1,2) < 3.0000000) ? 7.9999996M*V(1,2) + 182.99999M :
+ (V(1,2) < 3.5000000) ? 5.9999997M*V(1,2) + 188.99999M :
+ (V(1,2) < 4.0000000) ? 3.9999998M*V(1,2) + 195.99999M :
+ (V(1,2) < 4.5000000) ? 3.9999998M*V(1,2) + 195.99999M :
+ (V(1,2) < 5.0000000) ? 1.9999999M*V(1,2) + 204.99999M :
+ (V(1,2) < 10.0000000) ? 1.0000000M*V(1,2) + 209.99999M :
+ 1.0000000N*V(1,2) + 219.99998M
.ENDS
.SUBCKT PCIIW  4     300 400
*Connections    Input VCC VEE
* Diode Clamps
XVCC_OUT 6 300 300 6 VCC_OUT
XGND_OUT 6 400 6 400 GND_OUT
V5 6 5 
* Package Parasitics Max
ROSNB 5 1 100
ROPKG 1 4 .200
COPKG 4 400 2.00P
CCOMP 5 400 8.00P
LOPKG 5 1 15.00N
.ENDS
.SUBCKT GND_OUT  3    4    1   2
*                OUT+ OUT- IN+ IN-
B1 3 4 I= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + -292.99998M :
+ (V(1,2) < -1.0000000) ? 66.999997M*V(1,2) + 41.999998M :
+ (V(1,2) < -899.99996M) ? 119.99999M*V(1,2) + 94.999995M :
+ (V(1,2) < -799.99996M) ? 69.999997M*V(1,2) + 49.999998M :
+ (V(1,2) < -699.99997M) ? 35.999998M*V(1,2) + 22.799999M :
+ (V(1,2) < -599.99997M) ? 11.999999M*V(1,2) + 5.9999997M :
+ (V(1,2) < -499.99998M) ? 6.9999997M*V(1,2) + 2.9999999M :
+ (V(1,2) < -399.99998M) ? 3.9999998M*V(1,2) + 1.4999999M :
+ (V(1,2) < 0.0000000E+00) ? 250.00000U*V(1,2) + -6.6174449E-12 :
+ 1.0000000N*V(1,2) + 0.0000000E+00
.ENDS
*
.SUBCKT VCC_OUT 3    4    1   2
*               OUT+ OUT- IN+ IN-
B1 3 4 I= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + 292.99999M :
+ (V(1,2) < -1.0000000) ? -66.999997M*V(1,2) + -41.999998M :
+ (V(1,2) < -899.99996M) ? -119.99999M*V(1,2) + -94.999995M :
+ (V(1,2) < -799.99996M) ? -69.999997M*V(1,2) + -49.999998M :
+ (V(1,2) < -699.99997M) ? -35.999998M*V(1,2) + -22.799999M :
+ (V(1,2) < -599.99997M) ? -11.999999M*V(1,2) + -5.9999997M :
+ (V(1,2) < -499.99998M) ? -6.9999997M*V(1,2) + -2.9999999M :
+ (V(1,2) < -399.99998M) ? -3.9999998M*V(1,2) + -1.4999999M :
+ (V(1,2) < 0.0000000E+00) ? -250.00000U*V(1,2) + 6.6174449E-12 :
+ 1.0000000N*V(1,2) + 0.0000000E+00
.ENDS
*
.OPTION ACCT VSCALE=5
*INCLUDE FRAME.LIB
*ALIAS  V(100)=VINPUT
*ALIAS  V(500)=ENABLE
*ALIAS  V(1)=VTIN
*ALIAS  V(2)=VTOUT
.PRINT TRAN  V(100)  V(500)  V(1)  V(2) 
V2 500 0 5
V3 300 0 5
V4 400 0 0
X6 100 1 300 400 500 PCIOB
T1 1 0 2 0 ZO=65 TD=1.5N
X12 2 300 400 PCIIW
V1 100 0 PULSE 0 5 2N 2.5N 2.5N 50N 100N
.END
