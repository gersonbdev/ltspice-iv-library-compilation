*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Inc.
* Models developed and under copyright by:
* National Semiconductor, Inc.  

*/////////////////////////////////////////////////////////////////////
* Legal Notice: This material is intended for free software support.
* The file may be copied, and distributed; however, reselling the 
*  material is illegal

*////////////////////////////////////////////////////////////////////
* For ordering or technical information on these models, contact:
* National Semiconductor's Customer Response Center
*                 7:00 A.M.--7:00 P.M.  U.S. Central Time
*                                (800) 272-9959
* For Applications support, contact the Internet address:
*  amps-apps@galaxy.nsc.com

*//////////////////////////////////////////////////////////
*LMC6684B CMOS QUAD OP-AMP MACRO-MODEL
*//////////////////////////////////////////////////////////
*
* Connections:      Non-inverting input
*                   |   Inverting input
*                   |   |   Positive power supply
*                   |   |   |   Negative power supply
*                   |   |   |   |   Output
*                   |   |   |   |   |   Shutdown
*                   |   |   |   |   |   |
.SUBCKT LMC6684B/NS 1   2  99  50  28  33
* CAUTION:  SET .OPTIONS GMIN=1E-16 TO CORRECTLY MODEL INPUT BIAS CURRENT.
* Features:
* Operates from single supply
* Rail-to-rail output swing
* Low offset voltage (max) = 3mV@5V
* Slew rate = 1.2V/uS
* Gain-bandwidth product = 1.2 MHz 
* Amplifier shut-down
* Power is for one amplifier
*
* NOTE: - Model is for single device only and simulated.
*       - Noise is not modeled.
*       - Asymmetrical gain is not modeled.
*
CI1 1  50 2P
CI2 2  50 2P
* 1.4 Hz pole capacitor
C3  98 9  5.85N
* 2.95 MHz pole capacitor
C4  6  5  4.93P
* Drain-substrate capacitor
C6  50 4  10P
* 35 MHz pole capacitor
C7  98 11 4.54F
COUT 28 0 10P
CSD1 41 40 100P
DP1 1  99 DA
DP2 50 1  DX
DP3 2  99 DB
DP4 50 2  DX
D1  9  8  DX
D2  10 9  DX
D3  29 22 DX
D4  22 30 DX
D5  22 26 DX
D6  27 22 DX
D7  22 99 DX
D8  50 22 DX
D9  0  14 DX
D10 12 0  DX
D11 31 32 DX
EH  97 98 99    49 1.0
EN  0  96 0     50 1.0
* Input offset voltage -|
EOS 7  1  POLY(1) 16 49 3M 1
EP  97 0  99    0  1.0
E1  97 23 99    15 1.0
E2 18 7 32 97 1E-3
* Sourcing load +Vs current
F1  99 0  VA2   1
* Sinking load -Vs current
F2  0  50 VA3   1
F3  13 0  VA1   1
G1  98 9  5     6  0.1
G2  98 11 9     49 1U
G3  98 15 11    49 1U
* DC CMRR
G4  98 16 POLY(2) 1 49 2 49 0 3.54E-8 3.54E-8
G5  99 4  39 45 11.5U
G6  99 50 39 45 340U
* Load dependent pole
L1 19 28 40.4U
* CMR lead
L2  16 17 7.95M
M1  5  2  4     99 MPX
M2  6  18 4     99 MPX
M3 41 33 40 40 MN1
M4 45 41 39 39 MP2
M5 45 41 40 40 MN3 
R3  5  50 3.60K
R4  6  50 3.60K
R5  98 9  1E7
R8  42 44 25K
R9  44 50 25K
R12 98 11 1E6
R13 98 17 1K
* -Rout
R16 23 24 55
* +Rout
R17 23 25 55
* +Isc slope control
R18 15 20 1MEG
* -Isc slope control
R19 21 15 400K
R21 98 15 1E6
R22 19 28 900
R23 32 97 100K
R24 99 49 10MEG
R25 49 50 10MEG
R26 33 50 20MEG
R27 39 41 250K
S1 99 42 41 49 SX 
S2 22 36 41 49 SX
VA1 36 19 0V
VA2 14 13 0V
VA3 13 12 0V
V2  97 8  0.66V
V3  10 96 0.66V
V4  20 29 0.13V
V5  30 21 0.13V
V6  24 26 0.63V
V7  27 25 0.63V
V8 31 96 3.6V 
V9 39 49 1
V10 49 40 1
*
.MODEL DA D    (IS=250E-15)
.MODEL DB D    (IS=175E-15)
.MODEL DX D    (IS=100E-15)
.MODEL MPX PMOS (VTO=-.6 KP=7.0547E-4 GAMMA=1.1)
.MODEL MN1 NMOS (VTO=.6 KP=7.0547E-4 GAMMA=1.1)
.MODEL MP2 PMOS (VTO=0, KP=7.0547E-4)
.MODEL MN3 NMOS (VTO=0, KP=7.0547E-4)
.MODEL SX VSWITCH (RON=1, ROFF=1E+8, VON=0.01, VOFF=-0.01)
.ENDS
*
*$
