IBIS
*SPICE_NET
.TRAN .1N 120N
*INCLUDE IBIS1.LIB
.SUBCKT PCIIW  4     300 400
*Connections    Input VCC VEE
* Diode Clamps
XVCC_OUT 6 300 300 6 VCC_OUT
XGND_OUT 6 400 6 400 GND_OUT
V5 6 5 
* Package Parasitics Max
ROSNB 5 1 100
ROPKG 1 4 .200
COPKG 4 400 2.00P
CCOMP 5 400 8.00P
LOPKG 5 1 15.00N
.ENDS
.SUBCKT GND_OUT  3    4    1   2
*                OUT+ OUT- IN+ IN-
B1 3 4 I= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + -292.99998M :
+ (V(1,2) < -1.0000000) ? 66.999997M*V(1,2) + 41.999998M :
+ (V(1,2) < -899.99996M) ? 119.99999M*V(1,2) + 94.999995M :
+ (V(1,2) < -799.99996M) ? 69.999997M*V(1,2) + 49.999998M :
+ (V(1,2) < -699.99997M) ? 35.999998M*V(1,2) + 22.799999M :
+ (V(1,2) < -599.99997M) ? 11.999999M*V(1,2) + 5.9999997M :
+ (V(1,2) < -499.99998M) ? 6.9999997M*V(1,2) + 2.9999999M :
+ (V(1,2) < -399.99998M) ? 3.9999998M*V(1,2) + 1.4999999M :
+ (V(1,2) < 0.0000000E+00) ? 250.00000U*V(1,2) + -6.6174449E-12 :
+ 1.0000000N*V(1,2) + 0.0000000E+00
.ENDS
*
.SUBCKT VCC_OUT 3    4    1   2
*               OUT+ OUT- IN+ IN-
B1 3 4 I= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + 292.99999M :
+ (V(1,2) < -1.0000000) ? -66.999997M*V(1,2) + -41.999998M :
+ (V(1,2) < -899.99996M) ? -119.99999M*V(1,2) + -94.999995M :
+ (V(1,2) < -799.99996M) ? -69.999997M*V(1,2) + -49.999998M :
+ (V(1,2) < -699.99997M) ? -35.999998M*V(1,2) + -22.799999M :
+ (V(1,2) < -599.99997M) ? -11.999999M*V(1,2) + -5.9999997M :
+ (V(1,2) < -499.99998M) ? -6.9999997M*V(1,2) + -2.9999999M :
+ (V(1,2) < -399.99998M) ? -3.9999998M*V(1,2) + -1.4999999M :
+ (V(1,2) < 0.0000000E+00) ? -250.00000U*V(1,2) + 6.6174449E-12 :
+ 1.0000000N*V(1,2) + 0.0000000E+00
.ENDS
*
.SUBCKT PCIOW 100   4      300 400 500
*Connections    Input Output VCC VEE Enable
*Passed Parameters; Max
*dEFINE {RTF}=40K
*dEFINE {RTR}=40K
* Input Control
B1 820 0 V=V(100) & V(500)
B2 830 0 V= V(500) & ~V(100)
* Up and Down Ramps
B3 300 850 I= V(830) > 1.2   ? 0 : V(300,850) / 40K
B4 840 400 I= V(820) > 1.2 ? 0 : V(840,400) / 40K
C1 300 850 .01P
C2 840 400 .01P
S1 220 850 0 820 SMOD
S2 840 220 0 830 SMOD
.MODEL SMOD SW RON=.1M ROFF=1E15 VT=-1.2 VH=.1
G1 8 400 2 8 1
R1 6 400 1
G2 300 8 8 3 1
R2 300 6 1
* Pull-up/Pull-down structures; Min
XEPL_DN 2 400 8 840 EPWL_DNN
XEPL_UP 3 300 850 8 EPWL_UPN
* Diode Clamps
XVCC_OUT 6 300 300 6 VCC_OUT
XGND_OUT 6 400 6 400 GND_OUT
* Package Parasitics; Max
ROSNB 5 1 100
ROPKG 1 4 .200
COPKG 4 400 2.00P
CCOMP 5 400 8.00P
LOPKG 5 1 15.00N
* Voltage Sources for measuring currents
V5 6 5 
V6 8 6 
V7 220 8 
.ENDS
*Subcircuits for the IBIS1 Topology
.SUBCKT GND_OUT  3    4    1   2
*                OUT+ OUT- IN+ IN-
B1 3 4 I= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + -292.99998M :
+ (V(1,2) < -1.0000000) ? 66.999997M*V(1,2) + 41.999998M :
+ (V(1,2) < -899.99996M) ? 119.99999M*V(1,2) + 94.999995M :
+ (V(1,2) < -799.99996M) ? 69.999997M*V(1,2) + 49.999998M :
+ (V(1,2) < -699.99997M) ? 35.999998M*V(1,2) + 22.799999M :
+ (V(1,2) < -599.99997M) ? 11.999999M*V(1,2) + 5.9999997M :
+ (V(1,2) < -499.99998M) ? 6.9999997M*V(1,2) + 2.9999999M :
+ (V(1,2) < -399.99998M) ? 3.9999998M*V(1,2) + 1.4999999M :
+ (V(1,2) < 0.0000000E+00) ? 250.00000U*V(1,2) + -6.6174449E-12 :
+ 1.0000000N*V(1,2) + 0.0000000E+00
.ENDS
*
.SUBCKT VCC_OUT 3    4    1   2
*               OUT+ OUT- IN+ IN-
B1 3 4 I= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + 292.99999M :
+ (V(1,2) < -1.0000000) ? -66.999997M*V(1,2) + -41.999998M :
+ (V(1,2) < -899.99996M) ? -119.99999M*V(1,2) + -94.999995M :
+ (V(1,2) < -799.99996M) ? -69.999997M*V(1,2) + -49.999998M :
+ (V(1,2) < -699.99997M) ? -35.999998M*V(1,2) + -22.799999M :
+ (V(1,2) < -599.99997M) ? -11.999999M*V(1,2) + -5.9999997M :
+ (V(1,2) < -499.99998M) ? -6.9999997M*V(1,2) + -2.9999999M :
+ (V(1,2) < -399.99998M) ? -3.9999998M*V(1,2) + -1.4999999M :
+ (V(1,2) < 0.0000000E+00) ? -250.00000U*V(1,2) + 6.6174449E-12 :
+ 1.0000000N*V(1,2) + 0.0000000E+00
.ENDS
*
.SUBCKT EPWL_UPN 3    4    1   2
*                OUT+ OUT- IN+ IN-
B1 3 4 V= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + 55.000002M :
+ (V(1,2) < -4.0000000) ? -1.9999999M*V(1,2) + 44.999998M :
+ (V(1,2) < -3.0000000) ? -4.9999998M*V(1,2) + 32.999998M :
+ (V(1,2) < -2.0000000) ? -10.999999M*V(1,2) + 14.999999M :
+ (V(1,2) < -1.0000000) ? -14.999999M*V(1,2) + 6.9999997M :
+ (V(1,2) < 0.0000000E+00) ? -21.999999M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 499.99998M) ? -25.999999M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 1.0000000) ? -17.999999M*V(1,2) + -3.9999998M :
+ (V(1,2) < 1.5000000) ? -15.999999M*V(1,2) + -5.9999997M :
+ (V(1,2) < 2.0000000) ? -13.999999M*V(1,2) + -8.9999996M :
+ (V(1,2) < 2.5000000) ? -11.999999M*V(1,2) + -12.999999M :
+ (V(1,2) < 3.0000000) ? -9.9999995M*V(1,2) + -17.999999M :
+ (V(1,2) < 3.5000000) ? -5.9999997M*V(1,2) + -29.999999M :
+ (V(1,2) < 4.0000000) ? -3.9999998M*V(1,2) + -36.999998M :
+ (V(1,2) < 4.5000000) ? -1.9999999M*V(1,2) + -44.999998M :
+ (V(1,2) < 5.0000000) ? -1.9999999M*V(1,2) + -44.999998M :
+ (V(1,2) < 10.0000000) ? -400.00000U*V(1,2) + -52.999997M :
+ 1.0000000N*V(1,2) + -57.000007M
.ENDS
*
.SUBCKT EPWL_DNN  3    4    1   2
*                 OUT+ OUT- IN+ IN-
B1 3 4 V= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + -109.99999M :
+ (V(1,2) < -4.0000000) ? 1.9999999M*V(1,2) + -99.999995M :
+ (V(1,2) < -3.0000000) ? 4.9999998M*V(1,2) + -87.999996M :
+ (V(1,2) < -2.0000000) ? 10.999999M*V(1,2) + -69.999997M :
+ (V(1,2) < -1.0000000) ? 56.999997M*V(1,2) + 21.999999M :
+ (V(1,2) < 0.0000000E+00) ? 34.999998M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 499.99998M) ? 69.999997M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 1.0000000) ? 45.999998M*V(1,2) + 11.999999M :
+ (V(1,2) < 1.5000000) ? 35.999998M*V(1,2) + 21.999999M :
+ (V(1,2) < 2.0000000) ? 31.999998M*V(1,2) + 27.999999M :
+ (V(1,2) < 2.5000000) ? 15.999999M*V(1,2) + 59.999997M :
+ (V(1,2) < 3.0000000) ? 5.9999997M*V(1,2) + 84.999996M :
+ (V(1,2) < 3.5000000) ? 3.9999998M*V(1,2) + 90.999996M :
+ (V(1,2) < 4.0000000) ? 5.9999997M*V(1,2) + 83.999996M :
+ (V(1,2) < 4.5000000) ? 1.9999999M*V(1,2) + 99.999995M :
+ (V(1,2) < 5.0000000) ? 1.9999999M*V(1,2) + 99.999995M :
+ (V(1,2) < 10.0000000) ? 1.0000000M*V(1,2) + 105.00000M :
+ 1.0000000N*V(1,2) + 114.99998M
.ENDS
.SUBCKT BLINE#0 1 2 
*Interconnect Model for the Buried Microstrip PCI Speedway line
O1 1 0 2 0 LOSSY
.MODEL LOSSY LTRA rel=1.8 len=27.940MM
+ r=0 g=0
+ l=723NH/m
+ c=76PF/m 
* z0 = 97.535 Ohms 
* td = 7.4127Ns
* Total Delay = 207.11Ps
.ENDS
.SUBCKT BLINE#1 1 2 
*Interconnect Model for the Buried Microstrip PCI Speedway line
O1 1 0 2 0 LOSSY
.MODEL LOSSY LTRA rel=1.8 len=25.400MM
+ r=0 g=0
+ l=723NH/m
+ c=76PF/m 
* z0 = 97.535 Ohms 
* td = 7.4127Ns
* Total Delay = 188.28Ps
.ENDS
.SUBCKT BLINE#2 1 2 
*Interconnect Model for the Suface Microstrip Stub from the 
* PCI Speedway to the Load
O1 1 0 2 0 LOSSY
.MODEL LOSSY LTRA rel=1.8 len=40.640MM
+ r=0 g=0
+ l=523NH/m
+ c=76PF/m 
* z0 = 82.955 Ohms
* td = 6.3046Ns
* Total Delay = 256.22Ps
.ENDS
.SUBCKT BLINE#3 1 2 
*Interconnect Model for the Suface Microstrip Stub from the 
* PCI Speedway to the Load
O1 1 0 2 0 LOSSY
.MODEL LOSSY LTRA rel=1.8 len=38.100MM
+ r=0 g=0
+ l=523NH/m
+ c=76PF/m 
* z0 = 82.955 Ohms
* td = 6.3046Ns
* Total Delay = 240.21Ps
.ENDS
.OPTION ACCT VSCALE=7.5
*ALIAS  V(100)=VINPUT
*ALIAS  V(500)=ENABLE
*ALIAS  V(1)=VB
*ALIAS  V(14)=VA
*ALIAS  V(3)=VLOAD2
*ALIAS  V(17)=VLOAD10
.PRINT TRAN  V(100)  V(500)  V(1)  V(14) 
.PRINT TRAN  V(3)  V(17) 
X36 3 300 400 PCIIW
V1 100 0 PULSE 0 5 0 2.5N 2.5N 30N 60N
V2 500 0 5
V3 300 0 5.25
V4 400 0 0
X6 100 14 300 400 500 PCIOW
X16 100 1 300 400 500 PCIOW
C1 1 0 40PF
X32 9 300 400 PCIIW
X33 22 300 400 PCIIW
X34 23 300 400 PCIIW
X35 24 300 400 PCIIW
X37 6 300 400 PCIIW
X38 4 300 400 PCIIW
X39 8 300 400 PCIIW
C2 11 0 .5PF
C3 10 0 .5PF
C4 5 0 .5PF
C5 16 0 .5PF
C6 15 0 .5PF
C7 7 0 .5PF
C8 13 0 .5PF
C9 12 0 .5PF
C10 18 0 .5PF
X3 14 11 BLINE#0 
*{LENGTH=1.1 }
X97 11 7 BLINE#1 
*{LENGTH=1 }
X98 7 10 BLINE#1 
*{LENGTH=1 }
X99 10 13 BLINE#1 
*{LENGTH=1 }
X100 13 5 BLINE#1 
*{LENGTH=1 }
X101 5 12 BLINE#1 
*{LENGTH=1 }
X102 12 16 BLINE#1 
*{LENGTH=1 }
X103 16 18 BLINE#1 
*{LENGTH=1 }
X104 18 15 BLINE#1 
*{LENGTH=1 }
X105 3 11 BLINE#2 
*{LENGTH=1.6 }
X106 6 10 BLINE#3 
*{LENGTH=1.5 }
X107 4 5 BLINE#3 
*{LENGTH=1.5 }
X108 8 16 BLINE#3 
*{LENGTH=1.5 }
X109 17 15 BLINE#3 
*{LENGTH=1.5 }
X110 9 7 BLINE#3 
*{LENGTH=1.5 }
X111 22 13 BLINE#3 
*{LENGTH=1.5 }
X112 23 12 BLINE#3 
*{LENGTH=1.5 }
X113 24 18 BLINE#3 
*{LENGTH=1.5 }
X40 17 300 400 PCIIW
.END
