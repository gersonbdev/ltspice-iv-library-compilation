SCN3
.OPTIONS ACCT
*SPICE_NET
*INCLUDE DEVICE.LIB
.TRAN .05U 20U
.OPTIONS LIMPTS=20000 PIVTOL=1E-20
*ALIAS  V(2)=PHASE2
*ALIAS  V(1)=PHASE1
*ALIAS  V(14)=VOUT
.PRINT TRAN  V(2)  V(1)  V(14) 
X2 9 0 2 SWITCH 
X3 3 4 2 SWITCH 
X4 8 0 1 SWITCH 
X5 14 5 2 SWITCH 
X6 8 10 2 SWITCH 
X7 4 0 1 SWITCH 
X9 7 10 2 SWITCH 
X10 19 9 1 SWITCH 
C1 5 8 2P
C2 4 8 2P
C3 9 7 2P
X12 7 0 1 SWITCH 
X13 11 12 1 SWITCH 
X14 12 0 2 SWITCH 
X15 13 0 1 SWITCH 
X16 13 16 2 SWITCH 
E1 11 0 0 10 1K
C4 10 11 32P
C5 12 13 2P
E2 14 0 0 16 1K
C6 16 14 32P
E3 19 0 0 18 20K
R1 11 18 100K
R2 18 19 10K
V1 3 0 PULSE 0 2
V2 2 0 PULSE 0 1 0 0 0 0.8U 2U
V3 1 0 PULSE 0 1 1U 0 0 .8U 2U
R3 2 0 1K
R4 1 0 1K
X1 5 0 1 SWITCH 
.END