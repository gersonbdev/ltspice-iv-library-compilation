SCN13
.OPTIONS LIMPTS=1000
*SPICE_NET
*INCLUDE SCN.LIB
.SUBCKT SCNAMP64 2    3  6
*                - IN + OUT
*PARAMS ARE GAIN=80.000  FT=7.0000MEG IOS=1.0000P VOS=1.0000M IBIAS=3.0000P     
*GAIN IS IN db  
RIP 3 0 10MEG   
CIP 3 0 1.4PF   
IBN 2 0 3.0000P 
RIN 2 0 10MEG   
CIN 2 0 1.4PF   
VOFST 2 10 1.0000M      
RID 10 3 200K   
EA 11 0 10 3 1  
R1 11 12 5K     
R2 12 13 50K    
C1 12 0 1.8571P 
GA 0 14 0 13 135.00     
C2 13 14 385.71F
RO 14 0 75      
L 14 6 4.2857U  
RL 14 6 1000    
CL 6 0 3PF      
.ENDS   
.SUBCKT LT6450D 3 2 1 33 28 10 4 6 14 29 12 5 22 24 30 13 8 31 32 26 17
*Connections   INVA AGND HPA SA BPA LPA INVB HPB SB BPB LPB 
*Connections                    INVC HPC SC BPC LPC INVD HPD BPD LPD CLK
*Subcircuit for DIP package
X10 16 17 18 MUL#0  
*{K=1 } 
X11 28 17 20 MUL#0  
*{K=1 } 
X12 18 28 SINT#0  
*{K=62.5K } 
X13 20 10 SINT#0  
*{K=62.5K } 
X15 1 33 16 SUM2#0  
*{K1=1 K2=-1 }
X16 4 2 6 SCNAMP64
X17 7 17 9 MUL#0  
*{K=1 } 
X18 29 17 11 MUL#0  
*{K=1 } 
X19 9 29 SINT#0  
*{K=62.5K } 
X20 11 12 SINT#0  
*{K=62.5K } 
X21 6 14 7 SUM2#0  
*{K1=1 K2=-1 }
X22 5 2 22 SCNAMP64
X23 23 17 25 MUL#0  
*{K=1 } 
X24 30 17 27 MUL#0  
*{K=1 } 
X25 25 30 SINT#0  
*{K=62.5K } 
X26 27 13 SINT#0  
*{K=62.5K } 
X27 22 24 23 SUM2#0  
*{K1=1 K2=-1 }
X28 8 2 31 SCNAMP64
X29 31 17 34 MUL#0  
*{K=1 } 
X30 32 17 36 MUL#0  
*{K=1 } 
X31 34 32 SINT#0  
*{K=62.5K } 
X32 36 26 SINT#0  
*{K=62.5K } 
X5 3 2 1 SCNAMP64
.ENDS
*INCLUDE SYS.LIB
.SUBCKT MUL#0 1 2 3
RIN1 1 0 1E12
RIN2 2 0 1E12
ROUT 3 0 1E12
E1 3 0 POLY(2) 1 0 2 0 0 0 0 0 1.0000 
.ENDS
.SUBCKT SINT#0 1 2
*PARAMS ARE GAIN=62.500K
RIN 1 0 1E12
E1 3 0 0 1 62.500K
C1 2 4 1U IC=0
R1 3 4 1MEG
E2 2 0 0 4 1.0000MEG
.ENDS
.SUBCKT SUM2#0 1 2 3
RIN1 1 0 1E12
RIN2 2 0 1E12
ROUT 3 0 1E12
E1 3 0 POLY(2) 1 0 2 0 0 1.0000  -1.0000 
.ENDS
.AC DEC 100 1K 100K
*ALIAS  V(16)=VOUT
.PRINT AC  V(16)  VP(16) 
R12 12 14 46.95K
R14 15 20 10.5K
R15 16 20 39.42K
R16 17 20 13.19K
V2 14 0 AC 1
R17 1 5 10K
R18 3 5 70.3K
R19 2 5 16.3K
R20 1 20 17.9K
R21 2 20 69.7K
R22 4 5 27.46K
R23 7 5 6.9K
R24 7 8 10K
R25 6 8 81.5K
R26 4 8 14.72K
R27 8 25 93.93K
R28 12 10 11.81K
R29 12 25 38.25K
R30 12 11 10K
X2 12 0 11 0 25 10 8 7 0 6 4 5 2 0 3 1 20 17 16 15 9 LT6450D 
V1 9 0 2
.END