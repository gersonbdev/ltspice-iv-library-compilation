SCN11
.OPTIONS ITL5=0
*SPICE_NET
.TRAN .1M 50M
.OPTIONS ACCT LIMPTS=1000 PIVTOL=1E-20
*INCLUDE SCN.LIB
.SUBCKT SCNAMP60 2    3  6
*                - IN + OUT       
*PARAMS ARE GAIN=85.000  FT=2.0000MEG IOS=1.0000P VOS=1.0000M IBIAS=3.0000P     
*GAIN IS IN db  
RIP 3 0 10MEG   
CIP 3 0 1.4PF   
IBN 2 0 3.0000P 
RIN 2 0 10MEG   
CIN 2 0 1.4PF   
VOFST 2 10 1.0000M      
RID 10 3 200K   
EA 11 0 10 3 1  
R1 11 12 5K     
R2 12 13 50K    
C1 12 0 6.5000P 
GA 0 14 0 13 240.07     
C2 13 14 1.3500P
RO 14 0 75      
L 14 6 15.000U  
RL 14 6 1000    
CL 6 0 3PF      
.ENDS   
.SUBCKT LT60L100 4    15   3   5   2   1   17   19  20  10   11   18  16 
* Connections    INVA AGND HPA S1A BPA LPA INVB BPB LPB CLKA CLKB HPB S1B
*Gain = 100, SAB switch set low
X3 2 10 7 MUL#0  
*{K=1 } 
X1 14 10 9 MUL#0  
*{K=1 } 
X8 15 3 5 14 SUM3#0  
*{K1=-1 K2=1 K3=-1 } 
XE2 4 15 3 SCNAMP60
X9 9 2 SINT#0  
*{K=31.25K } 
X10 7 1 SINT#0  
*{K=31.25K } 
*
X12 6 11 13 MUL#0  
*{K=1 } 
X13 19 11 22 MUL#0  
*{K=1 } 
XE3 17 15 18 SCNAMP60
X15 13 19 SINT#0  
*{K=31.25K } 
X16 22 20 SINT#0  
*{K=31.25K } 
X14 15 18 16 6 SUM3#0  
*{K1=-1 K2=1 K3=-1 } 
.ENDS
*INCLUDE SYS.LIB
.SUBCKT MUL#0 1 2 3
RIN1 1 0 1E12
RIN2 2 0 1E12
ROUT 3 0 1E12
E1 3 0 POLY(2) 1 0 2 0 0 0 0 0 1.0000 
.ENDS
.SUBCKT SUM3#0 1 2 3 4
* 3 PORT SUMMER
RIN1 1 0 1E12
RIN2 2 0 1E12
RIN3 3 0 1E12
ROUT 4 0 1E12
E1 4 0 POLY(3) 1 0 2 0 3 0 0 -1.0000  1.0000  -1.0000 
.ENDS
.SUBCKT SINT#0 1 2
*PARAMS ARE GAIN=31.250K
RIN 1 0 1E12
E1 3 0 0 1 31.250K
C1 2 4 1U IC=0
R1 3 4 1MEG
E2 2 0 0 4 1.0000MEG
.ENDS
*INCLUDE LIN.LIB 
.SUBCKT UA741 2    3  6   7   4
*             - IN + OUT VCC VEE
RP 4 7 10K
RXX 4 0 10MEG
*
IBP 3 0 80NA
RIP 3 0 10MEG
CIP 3 0 1.4PF
IBN 2 0 100NA
RIN 2 0 10MEG
CIN 2 0 1.4PF
VOFST 2 10 1MV
RID 10 3 200K
EA 11 0 10 3 1
R1 11 12 5K
R2 12 13 50K
C1 12 0 13PF
GA 0 14 0 13 2700
C2 13 14 2.7PF
RO 14 0 75
L 14 6 30UHY
RL 14 6 1000
CL 6 0 3PF
.ENDS
*ALIAS  V(4)=VSIG
*ALIAS  V(15)=VOUT
*ALIAS  V(9)=VL1
*ALIAS  V(12)=VL2
*ALIAS  V(13)=VCLK
.PRINT AC  V(15)  VP(15)  V(9)  VP(9) 
.PRINT AC  V(12)  VP(12) 
.PRINT TRAN  V(4)  V(15)  V(9)  V(12) 
.PRINT TRAN  V(13) 
R1 1 4 1K
R2 4 0 1K
V2 5 0 SFFM 0 1 900 5 2700
R3 5 4 1K
R4 4 6 155.93K
R5 6 7 5K
R6 6 8 152K
R7 6 9 5.27K
R8 9 10 10.74K
R9 7 10 13.2K
R10 10 14 5.26K
R11 10 11 151.8K
R12 10 12 5K
X2 17 0 15 18 19 UA741
V4 19 0 -15
V5 18 0 15
R13 14 17 5K
R14 17 15 37.3K
R15 12 17 6.11K
V6 13 0 SIN .04 .4 10
*SET TO 1 FOR 500KHZ, GAIN = 100 (100K,50)=.4 
C1 6 9 12P
C2 10 12 20P
X5 6 0 7 0 8 9 10 11 12 13 13 14 0 LT60L100 
V1 1 0 SFFM 0 1 100 5 300
.END