IBIS3
.SUBCKT NAND2 1 2 3
B1 3 0 V= ~(V(1) & V(2))
.ENDS
.SUBCKT AND2X 1 2 3
B1 3 0 V= (V(1) & ~V(2))
.ENDS
.SUBCKT DRVR 1  2  3   4
*            IN VCC VEE OUT
RC 4 3 1MEG
CC 4 3 1P
B1 0 4 I= V(1) > 1.2 ? V(2,4)/200 : V(3,4)/150
.ENDS
*SPICE_NET
.TRAN .1N 50N
.OPTIONS ACCT 
*ALIAS  V(14)=VOUT
*ALIAS  V(8)=VENABLE
*ALIAS  V(10)=VIN
*ALIAS  V(2)=VGUP
*ALIAS  V(5)=VGDN
*ALIAS  I(V5)=IDIE
*ALIAS  V(16)=VLGDN
*ALIAS  V(1)=VLGUP
*ALIAS  I(V6)=ICC
*ALIAS  V(7)=VDIE
.PRINT TRAN  V(14)  V(8)  V(10)  V(2) 
.PRINT TRAN  V(5)  I(V5) V(16)  V(1) 
.PRINT TRAN  I(V6) V(7) 
V2 8 0 PULSE 0 5 0 0 0 5N 10N
M1 7 5 9 9 NFET
.MODEL NFET NMOS CGDO=12N KP=.03 VTO=2.2
D1 7 4 DIODE
.MODEL DIODE D
D2 9 7 DIODE
C1 11 9 5.64P
L1 11 13 32.75N
R1 11 13 100
R2 13 14 .277
C2 14 9 1.36P
V3 9 0 
V4 6 0 5
V5 7 11 
X12 1 4 9 2 DRVR
X13 16 4 9 5 DRVR
X16 8 10 16 AND2X
V6 6 4 
R6 4 7 33K
R7 7 9 33K
M2 7 2 4 4 PFET
.MODEL PFET PMOS CGDO=12N KP=.015 VTO=-2.2
X17 10 8 1 NAND2
V1 10 0 PULSE 0 5 0 0 0 10N 20N
.END
