IBIS
*SPICE_NET
.TRAN .1N 150N
*INCLUDE IBIS1.LIB
.OPTION ACCT VSCALE=5
*INCLUDE FRAME.LIB
*ALIAS  V(100)=VINPUT
*ALIAS  V(500)=ENABLE
*ALIAS  V(1)=VTIN
*ALIAS  V(2)=VTOUT
.PRINT TRAN  V(100)  V(500)  V(1)  V(2) 
V2 500 0 5
V3 300 0 5
V4 400 0 0
X6 100 1 300 400 500 PCIOB
T1 1 0 2 0 ZO=65 TD=1.5N
X12 2 300 400 PCIIW
V1 100 0 PULSE 0 5 2N 2.5N 2.5N 50N 100N
.END
