SCN11
.OPTIONS ITL5=0
*SPICE_NET
.TRAN .1M 50M
.OPTIONS ACCT LIMPTS=1000 PIVTOL=1E-20
*INCLUDE SCN.LIB
*INCLUDE LIN.LIB 
*ALIAS  V(4)=VSIG
*ALIAS  V(15)=VOUT
*ALIAS  V(9)=VL1
*ALIAS  V(12)=VL2
*ALIAS  V(13)=VCLK
.PRINT AC  V(15)  VP(15)  V(9)  VP(9) 
.PRINT AC  V(12)  VP(12) 
.PRINT TRAN  V(4)  V(15)  V(9)  V(12) 
.PRINT TRAN  V(13) 
R1 1 4 1K
R2 4 0 1K
V2 5 0 SFFM 0 1 900 5 2700
R3 5 4 1K
R4 4 6 155.93K
R5 6 7 5K
R6 6 8 152K
R7 6 9 5.27K
R8 9 10 10.74K
R9 7 10 13.2K
R10 10 14 5.26K
R11 10 11 151.8K
R12 10 12 5K
X2 17 0 15 18 19 UA741
V4 19 0 -15
V5 18 0 15
R13 14 17 5K
R14 17 15 37.3K
R15 12 17 6.11K
V6 13 0 SIN .04 .4 10
*SET TO 1 FOR 500KHZ, GAIN = 100 (100K,50)=.4 
C1 6 9 12P
C2 10 12 20P
X5 6 0 7 0 8 9 10 11 12 13 13 14 0 LT60L100 
V1 1 0 SFFM 0 1 100 5 300
.END