IBIS
*SPICE_NET
.TRAN .1N 120N
*INCLUDE IBIS1.LIB
.SUBCKT PCIOW 100   4      300 400 500
*Connections    Input Output VCC VEE Enable
*Passed Parameters; Max
*dEFINE {RTF}=40K
*dEFINE {RTR}=40K
* Input Control
B1 820 0 V=V(100) & V(500)
B2 830 0 V= V(500) & ~V(100)
* Up and Down Ramps
B3 300 850 I= V(830) > 1.2   ? 0 : V(300,850) / 40K
B4 840 400 I= V(820) > 1.2 ? 0 : V(840,400) / 40K
C1 300 850 .01P
C2 840 400 .01P
S1 220 850 0 820 SMOD
S2 840 220 0 830 SMOD
.MODEL SMOD SW RON=.1M ROFF=1E15 VT=-1.2 VH=.1
G1 8 400 2 8 1
R1 6 400 1
G2 300 8 8 3 1
R2 300 6 1
* Pull-up/Pull-down structures; Min
XEPL_DN 2 400 8 840 EPWL_DNN
XEPL_UP 3 300 850 8 EPWL_UPN
* Diode Clamps
XVCC_OUT 6 300 300 6 VCC_OUT
XGND_OUT 6 400 6 400 GND_OUT
* Package Parasitics; Max
ROSNB 5 1 100
ROPKG 1 4 .200
COPKG 4 400 2.00P
CCOMP 5 400 8.00P
LOPKG 5 1 15.00N
* Voltage Sources for measuring currents
V5 6 5 
V6 8 6 
V7 220 8 
.ENDS
*Subcircuits for the IBIS1 Topology
.SUBCKT GND_OUT  3    4    1   2
*                OUT+ OUT- IN+ IN-
B1 3 4 I= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + -292.99998M :
+ (V(1,2) < -1.0000000) ? 66.999997M*V(1,2) + 41.999998M :
+ (V(1,2) < -899.99996M) ? 119.99999M*V(1,2) + 94.999995M :
+ (V(1,2) < -799.99996M) ? 69.999997M*V(1,2) + 49.999998M :
+ (V(1,2) < -699.99997M) ? 35.999998M*V(1,2) + 22.799999M :
+ (V(1,2) < -599.99997M) ? 11.999999M*V(1,2) + 5.9999997M :
+ (V(1,2) < -499.99998M) ? 6.9999997M*V(1,2) + 2.9999999M :
+ (V(1,2) < -399.99998M) ? 3.9999998M*V(1,2) + 1.4999999M :
+ (V(1,2) < 0.0000000E+00) ? 250.00000U*V(1,2) + -6.6174449E-12 :
+ 1.0000000N*V(1,2) + 0.0000000E+00
.ENDS
*
.SUBCKT VCC_OUT 3    4    1   2
*               OUT+ OUT- IN+ IN-
B1 3 4 I= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + 292.99999M :
+ (V(1,2) < -1.0000000) ? -66.999997M*V(1,2) + -41.999998M :
+ (V(1,2) < -899.99996M) ? -119.99999M*V(1,2) + -94.999995M :
+ (V(1,2) < -799.99996M) ? -69.999997M*V(1,2) + -49.999998M :
+ (V(1,2) < -699.99997M) ? -35.999998M*V(1,2) + -22.799999M :
+ (V(1,2) < -599.99997M) ? -11.999999M*V(1,2) + -5.9999997M :
+ (V(1,2) < -499.99998M) ? -6.9999997M*V(1,2) + -2.9999999M :
+ (V(1,2) < -399.99998M) ? -3.9999998M*V(1,2) + -1.4999999M :
+ (V(1,2) < 0.0000000E+00) ? -250.00000U*V(1,2) + 6.6174449E-12 :
+ 1.0000000N*V(1,2) + 0.0000000E+00
.ENDS
*
.SUBCKT EPWL_UPN 3    4    1   2
*                OUT+ OUT- IN+ IN-
B1 3 4 V= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + 55.000002M :
+ (V(1,2) < -4.0000000) ? -1.9999999M*V(1,2) + 44.999998M :
+ (V(1,2) < -3.0000000) ? -4.9999998M*V(1,2) + 32.999998M :
+ (V(1,2) < -2.0000000) ? -10.999999M*V(1,2) + 14.999999M :
+ (V(1,2) < -1.0000000) ? -14.999999M*V(1,2) + 6.9999997M :
+ (V(1,2) < 0.0000000E+00) ? -21.999999M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 499.99998M) ? -25.999999M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 1.0000000) ? -17.999999M*V(1,2) + -3.9999998M :
+ (V(1,2) < 1.5000000) ? -15.999999M*V(1,2) + -5.9999997M :
+ (V(1,2) < 2.0000000) ? -13.999999M*V(1,2) + -8.9999996M :
+ (V(1,2) < 2.5000000) ? -11.999999M*V(1,2) + -12.999999M :
+ (V(1,2) < 3.0000000) ? -9.9999995M*V(1,2) + -17.999999M :
+ (V(1,2) < 3.5000000) ? -5.9999997M*V(1,2) + -29.999999M :
+ (V(1,2) < 4.0000000) ? -3.9999998M*V(1,2) + -36.999998M :
+ (V(1,2) < 4.5000000) ? -1.9999999M*V(1,2) + -44.999998M :
+ (V(1,2) < 5.0000000) ? -1.9999999M*V(1,2) + -44.999998M :
+ (V(1,2) < 10.0000000) ? -400.00000U*V(1,2) + -52.999997M :
+ 1.0000000N*V(1,2) + -57.000007M
.ENDS
*
.SUBCKT EPWL_DNN  3    4    1   2
*                 OUT+ OUT- IN+ IN-
B1 3 4 V= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + -109.99999M :
+ (V(1,2) < -4.0000000) ? 1.9999999M*V(1,2) + -99.999995M :
+ (V(1,2) < -3.0000000) ? 4.9999998M*V(1,2) + -87.999996M :
+ (V(1,2) < -2.0000000) ? 10.999999M*V(1,2) + -69.999997M :
+ (V(1,2) < -1.0000000) ? 56.999997M*V(1,2) + 21.999999M :
+ (V(1,2) < 0.0000000E+00) ? 34.999998M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 499.99998M) ? 69.999997M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 1.0000000) ? 45.999998M*V(1,2) + 11.999999M :
+ (V(1,2) < 1.5000000) ? 35.999998M*V(1,2) + 21.999999M :
+ (V(1,2) < 2.0000000) ? 31.999998M*V(1,2) + 27.999999M :
+ (V(1,2) < 2.5000000) ? 15.999999M*V(1,2) + 59.999997M :
+ (V(1,2) < 3.0000000) ? 5.9999997M*V(1,2) + 84.999996M :
+ (V(1,2) < 3.5000000) ? 3.9999998M*V(1,2) + 90.999996M :
+ (V(1,2) < 4.0000000) ? 5.9999997M*V(1,2) + 83.999996M :
+ (V(1,2) < 4.5000000) ? 1.9999999M*V(1,2) + 99.999995M :
+ (V(1,2) < 5.0000000) ? 1.9999999M*V(1,2) + 99.999995M :
+ (V(1,2) < 10.0000000) ? 1.0000000M*V(1,2) + 105.00000M :
+ 1.0000000N*V(1,2) + 114.99998M
.ENDS
.OPTION ACCT VSCALE=5
*INCLUDE FRAME.LIB
*ALIAS  V(100)=VINPUT
*ALIAS  V(500)=ENABLE
*ALIAS  V(7)=VOUT
.PRINT TRAN  V(100)  V(500)  V(7) 
V2 500 0 5
V3 300 0 5
V4 400 0 0
X6 100 7 300 400 500 PCIOW
C1 7 0 50PF
V1 100 0 PULSE 0 5 0 2.5N 2.5N 27.44N 59.88N
.END
