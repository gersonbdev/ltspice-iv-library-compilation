IBIS2
.OPTIONS VSCALE=5
.SUBCKT INV 1 2
* LOAD SET TO MAKE 0 AND 1 WITHIN 1PPM OF DESIRED VALUE
RIN1 1 0 3E8
E1 2 0  1 0 1 -1
.ENDS
.SUBCKT NSWITCH 1 2 3
R1 1 2 3E13
G1 1 2 POLY(2) 1 2 3 0 0 0 0 0 6.67M
* 150 OHM ON, 3E13 OFF
.ENDS
.SUBCKT SWITCH 1 2 3
R1 1 2 3E13
G1 1 2 POLY(2) 1 2 3 0 0 0 0 0 5M
* 200 OHM ON, 3E13 OFF
.ENDS
*SPICE_NET
.TRAN .1N 50N
.OPTIONS ACCT
*ALIAS  V(15)=VOUT
*ALIAS  V(13)=VENABLE
*ALIAS  V(16)=VIN
*ALIAS  V(1)=VGUP
*ALIAS  V(4)=VGDN
*ALIAS  I(V5)=IDIE
.PRINT TRAN  V(15)  V(13)  V(16)  V(1) 
.PRINT TRAN  V(4)  I(V5)
X3 1 5 8 NSWITCH
X4 9 4 6 SWITCH
X5 4 5 3 NSWITCH
X6 6 3 INV
X7 13 8 16 SWITCH
X8 13 6 7 SWITCH
X9 16 7 INV
V1 16 0 PULSE 0 1 0 0 0 10N 20N
V2 13 0 PULSE 0 1 0 0 0 5N 10N
M2 17 4 5 5 NFET
.MODEL NFET NMOS CGDO=12N KP=.03 VTO=2.2
M3 17 1 9 9 PFET
.MODEL PFET PMOS CGDO=12N KP=.015 VTO=-2.2
X10 9 1 2 SWITCH
D1 17 9 DIODE
.MODEL DIODE D
D2 5 17 DIODE
C1 10 5 5.64P
L1 10 14 32.75N
R1 10 14 100
R2 14 15 .277
C2 15 5 1.36P
V3 5 0 
V4 9 0 5
V5 17 10 
R3 9 17 33K
R4 17 5 33K
C3 4 5 1P
C4 9 1 1P
X1 8 2 INV
.END
