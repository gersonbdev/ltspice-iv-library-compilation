SCN9
*SPICE_NET
*INCLUDE SCN.LIB
.SUBCKT SCNAMP60 2    3  6
*                - IN + OUT       
*PARAMS ARE GAIN=85.000  FT=2.0000MEG IOS=1.0000P VOS=1.0000M IBIAS=3.0000P     
*GAIN IS IN db  
RIP 3 0 10MEG   
CIP 3 0 1.4PF   
IBN 2 0 3.0000P 
RIN 2 0 10MEG   
CIN 2 0 1.4PF   
VOFST 2 10 1.0000M      
RID 10 3 200K   
EA 11 0 10 3 1  
R1 11 12 5K     
R2 12 13 50K    
C1 12 0 6.5000P 
GA 0 14 0 13 240.07     
C2 13 14 1.3500P
RO 14 0 75      
L 14 6 15.000U  
RL 14 6 1000    
CL 6 0 3PF      
.ENDS   
.SUBCKT LT60L100 4    15   3   5   2   1   17   19  20  10   11   18  16 
* Connections    INVA AGND HPA S1A BPA LPA INVB BPB LPB CLKA CLKB HPB S1B
*Gain = 100, SAB switch set low
X3 2 10 7 MUL#0  
*{K=1 } 
X1 14 10 9 MUL#0  
*{K=1 } 
X8 15 3 5 14 SUM3#0  
*{K1=-1 K2=1 K3=-1 } 
XE2 4 15 3 SCNAMP60
X9 9 2 SINT#0  
*{K=31.25K } 
X10 7 1 SINT#0  
*{K=31.25K } 
*
X12 6 11 13 MUL#0  
*{K=1 } 
X13 19 11 22 MUL#0  
*{K=1 } 
XE3 17 15 18 SCNAMP60
X15 13 19 SINT#0  
*{K=31.25K } 
X16 22 20 SINT#0  
*{K=31.25K } 
X14 15 18 16 6 SUM3#0  
*{K1=-1 K2=1 K3=-1 } 
.ENDS
*INCLUDE SYS.LIB
.SUBCKT MUL#0 1 2 3
RIN1 1 0 1E12
RIN2 2 0 1E12
ROUT 3 0 1E12
E1 3 0 POLY(2) 1 0 2 0 0 0 0 0 1.0000 
.ENDS
.SUBCKT SUM3#0 1 2 3 4
* 3 PORT SUMMER
RIN1 1 0 1E12
RIN2 2 0 1E12
RIN3 3 0 1E12
ROUT 4 0 1E12
E1 4 0 POLY(3) 1 0 2 0 3 0 0 -1.0000  1.0000  -1.0000 
.ENDS
.SUBCKT SINT#0 1 2
*PARAMS ARE GAIN=31.250K
RIN 1 0 1E12
E1 3 0 0 1 31.250K
C1 2 4 1U IC=0
R1 3 4 1MEG
E2 2 0 0 4 1.0000MEG
.ENDS
*INCLUDE NONLIN.LIB
.SUBCKT UA741 2    3  6   7  4
*             - IN + OUT VCC VEE
*
QNI1 10 2 13 QNI1
QNI2 12 3 13 QNI2
.MODEL QNI1 NPN(NF=1.5 BF=111 IS=8E-16 CJE=3PF)
.MODEL QNI2 NPN(NF=1.5 BF=144 IS=8.3E-16 CJE=3PF)
Q3 13 14 4 QN741
IEE 4 14 185NA
CCM 13 4 2.5PF
RCM 13 4 10MEG
RC1 11 10 1K
RC2 11 12 1K
CHF 10 12 55PF
D1 7 11 D741
RP 7 4 10K
GA 0 15 12 10 .9MMHO
GCM 0 15 13 0 6.3NMHOS
R2 15 0 100K
D2 15 0 D741 OFF
D3 0 15 D741 OFF
C2 15 16 30PF
GB 16 0 15 0 12.5
RO2 16 0 1000
D4 16 17 D741P OFF
EP 17 0 7 0 -1.8 1
D5 18 16 D741P OFF
EN 0 18 0 4 -2.3 1
.MODEL D741P D(RS=1M)
D6 19 16 D741
D7 16 20 D741
IRO 20 19 170UA
RR0 16 21 1MEG
Q4 7 19 21 QNO
Q5 4 20 21 QPO
.MODEL QNO NPN(BF=150 CJC=3P IS=1E-14)
.MODEL QPO PNP(BF=150 CJC=3P IS=1E-14)
L1 21 6 30UHY
RL1 21 6 1K
.MODEL D741 D(CJO=3PF)
.MODEL QN741 NPN
.ENDS
.AC LIN 200 1.5K 2.5K
.OPTIONS ACCT PIVTOL=1E-20 LIMPTS=1000
*ALIAS  V(13)=VOUT
*ALIAS  V(1)=VL1
*ALIAS  V(6)=VL2
.PRINT AC  V(13)  VP(13)  V(1)  VP(1) 
.PRINT AC  V(6)  VP(6) 
.PRINT TRAN  V(13)  V(1)  V(6) 
R21 3 2 5K
R31 3 5 152K
R41 3 1 5.27K
RL1 1 7 10.74K
V1 4 0 PULSE 0 1 AC 1
RH1 2 7 13.2K
R22 7 9 5.26K
R32 7 10 151.8K
R42 7 6 5K
X2 15 0 13 11 12 UA741
V2 12 0 -15
V3 11 0 15
RH2 9 15 5K
RG 15 13 37.3K
RL2 6 15 6.11K
VCLK 14 0 .4
*SET TO .4 FOR 2KHz NATURAL FREQUENCY 
*SET TO 1 FOR 500KHZ, GAIN = 100
*SET TO 4 FOR 20KHz NATURAL FREQUENCY 
C1 3 1 12P
C2 7 6 20P
X3 3 0 2 0 5 1 7 10 6 14 14 9 0 LT60L100 
R11 4 3 155.93K
.END