scn5
*DEFINE /SCNCAP=2P
*SPICE_NET
*INCLUDE SYS.LIB
.SUBCKT MUL#0 1 2 3
RIN1 1 0 1E12
RIN2 2 0 1E12
ROUT 3 0 1E12
E1 3 0 POLY(2) 1 0 2 0 0 0 0 0 1.0000 
.ENDS
.SUBCKT SINT#0 1 2
*PARAMS ARE GAIN=31.250K
RIN 1 0 1E12
E1 3 0 0 1 31.250K
C1 2 4 1U IC=0
R1 3 4 1MEG
E2 2 0 0 4 1.0000MEG
.ENDS
.SUBCKT SUM3#0 1 2 3 4
* 3 PORT SUMMER
RIN1 1 0 1E12
RIN2 2 0 1E12
RIN3 3 0 1E12
ROUT 4 0 1E12
E1 4 0 POLY(3) 1 0 2 0 3 0 0 -1.0000  1.0000  -1.0000 
.ENDS
*INCLUDE SCN.LIB
*INCLUDE LIN.LIB
.SUBCKT OP1#0 2    3  6   7   4
*              - IN + OUT VCC VEE
*PARAMS ARE GAIN=85.000  FT=2.0000MEG IOS=1.0000P VOS=1.0000M IBIAS=3.0000P
*GAIN IS IN db
RP 4 7 10K
RXX 4 0 10MEG
*
IBP 3 0 2.0000P
RIP 3 0 10MEG
CIP 3 0 1.4PF
IBN 2 0 3.0000P
RIN 2 0 10MEG
CIN 2 0 1.4PF
VOFST 2 10 1.0000M
RID 10 3 200K
EA 11 0 10 3 1
R1 11 12 5K
R2 12 13 50K
C1 12 0 6.5000P
GA 0 14 0 13 240.07 
C2 13 14 1.3500P
RO 14 0 75
L 14 6 15.000U
RL 14 6 1000
CL 6 0 3PF
.ENDS
.SUBCKT OP1#1 2    3  6   7   4
*              - IN + OUT VCC VEE
*PARAMS ARE GAIN=80.000  FT=2.0000MEG IOS=1.0000P VOS=1.0000M IBIAS=3.0000P
*GAIN IS IN db
RP 4 7 10K
RXX 4 0 10MEG
*
IBP 3 0 2.0000P
RIP 3 0 10MEG
CIP 3 0 1.4PF
IBN 2 0 3.0000P
RIN 2 0 10MEG
CIN 2 0 1.4PF
VOFST 2 10 1.0000M
RID 10 3 200K
EA 11 0 10 3 1
R1 11 12 5K
R2 12 13 50K
C1 12 0 6.5000P
GA 0 14 0 13 135.00 
C2 13 14 1.3500P
RO 14 0 75
L 14 6 15.000U
RL 14 6 1000
CL 6 0 3PF
.ENDS
.SUBCKT OP1#2 2    3  6   7   4
*              - IN + OUT VCC VEE
*PARAMS ARE GAIN=80.000  FT=7.0000MEG IOS=1.0000P VOS=1.0000M IBIAS=3.0000P
*GAIN IS IN db
RP 4 7 10K
RXX 4 0 10MEG
*
IBP 3 0 2.0000P
RIP 3 0 10MEG
CIP 3 0 1.4PF
IBN 2 0 3.0000P
RIN 2 0 10MEG
CIN 2 0 1.4PF
VOFST 2 10 1.0000M
RID 10 3 200K
EA 11 0 10 3 1
R1 11 12 5K
R2 12 13 50K
C1 12 0 1.8571P
GA 0 14 0 13 135.00 
C2 13 14 385.71F
RO 14 0 75
L 14 6 4.2857U
RL 14 6 1000
CL 6 0 3PF
.ENDS
.SUBCKT OP1#3 2    3  6   7   4
*              - IN + OUT VCC VEE
*PARAMS ARE GAIN=83.000  FT=2.5000MEG IOS=1.0000P VOS=5.0000M IBIAS=10.0000P
*GAIN IS IN db
RP 4 7 10K
RXX 4 0 10MEG
*
IBP 3 0 9.0000P
RIP 3 0 10MEG
CIP 3 0 1.4PF
IBN 2 0 10.0000P
RIN 2 0 10MEG
CIN 2 0 1.4PF
VOFST 2 10 5.0000M
RID 10 3 200K
EA 11 0 10 3 1
R1 11 12 5K
R2 12 13 50K
C1 12 0 5.2000P
GA 0 14 0 13 190.69 
C2 13 14 1.0800P
RO 14 0 75
L 14 6 12.000U
RL 14 6 1000
CL 6 0 3PF
.ENDS
.SUBCKT OP1#4 2    3  6   7   4
*              - IN + OUT VCC VEE
*PARAMS ARE GAIN=80.000  FT=2.5000MEG IOS=1.0000P VOS=5.0000M IBIAS=10.0000P
*GAIN IS IN db
RP 4 7 10K
RXX 4 0 10MEG
*
IBP 3 0 9.0000P
RIP 3 0 10MEG
CIP 3 0 1.4PF
IBN 2 0 10.0000P
RIN 2 0 10MEG
CIN 2 0 1.4PF
VOFST 2 10 5.0000M
RID 10 3 200K
EA 11 0 10 3 1
R1 11 12 5K
R2 12 13 50K
C1 12 0 5.2000P
GA 0 14 0 13 135.00 
C2 13 14 1.0800P
RO 14 0 75
L 14 6 12.000U
RL 14 6 1000
CL 6 0 3PF
.ENDS
.SUBCKT OPAMP#0 2    3  6   7   4
*             - IN + OUT VCC VEE
*PARAMS ARE GAIN=28.000K FT=2.5000MEG IOS=1.0000P VOS=0.0000E0 IBIAS=1.0000P
RP 4 7 10K
RXX 4 0 10MEG
*
IBP 3 0 0.0000E0
RIP 3 0 10MEG
CIP 3 0 1.4PF
IBN 2 0 1.0000P
RIN 2 0 10MEG
CIN 2 0 1.4PF
VOFST 2 10 0.0000E0
RID 10 3 200K
EA 11 0 10 3 1
R1 11 12 5K
R2 12 13 50K
C1 12 0 5.2000P
GA 0 14 0 13 378.00 
C2 13 14 1.0800P
RO 14 0 75
L 14 6 12.000U
RL 14 6 1000
CL 6 0 3PF
.ENDS
X12 6 11 13 MUL#0  
*{K=1 } 
X13 19 11 22 MUL#0  
*{K=1 } 
X15 13 19 SINT#0  
*{K=31.25K } 
X16 22 20 SINT#0  
*{K=31.25K } 
X18 20 4 16 7 SUM3#0  
*{K1=-1 K2=1 K3=-1 } 
X19 7 8 9 MUL#0  
*{K=1 } 
X20 19 8 14 MUL#0  
*{K=1 } 
X21 9 19 SINT#0  
*{K=31.25K } 
X22 14 20 SINT#0  
*{K=31.25K } 
X14 24 1 16 6 SUM3#0  
*{K1=-1 K2=1 K3=-1 } 
*
X17 2 3 1 7 4 OP1#0 
*{IBIAS=3P IOS=1P VOS=1M GAIN=85 FT=2MEG}
*LTC1060
X17 2 3 1 7 4 OP1#1 
*{IBIAS=3P IOS=1P VOS=1M GAIN=80 FT=2MEG}
*LTC1059
X17 2 3 1 7 4 OP1#2 
*{IBIAS=3P IOS=1P VOS=1M GAIN=80 FT=7MEG}
*LTC1064
X17 2 3 1 7 4 OP1#3 
*{IBIAS=10P IOS=1P VOS=5M GAIN=83 FT=2.5MEG}
*MF10
X17 2 3 1 7 4 OP1#4 
*{IBIAS=10P IOS=1P VOS=5M GAIN=80 FT=2.5MEG}
*MF5
X17 2 3 1 7 4 OPAMP#0 
*{IBIAS=1P IOS=1P VOS=0M GAIN=28000 FT=2.5MEG}
*TEST
.END