SCN2
*SPICE_NET
*INCLUDE SCN.LIB
.SUBCKT CRES#0 1 2
R1 1 2 500.00 
.ENDS

.SUBCKT NSTR#0 1 2
*NEGATIVE STORISTER I = 1E9 * (- C * Z^-1/2)
E1 3 0 1 2 1
T1 3 0 4 0 Z0=1000 TD=1.0000U
RT 4 0 1000
G1 1 2 0 4 2.0000M
.ENDS
.SUBCKT ZINT#0 1 2 3 4 
* 2 PHASE INT, 1 3 ARE ODD IN->OUT; 2,4 ARE EVEN
R1 1 3 31.250 
R2 2 4 31.250 

E13 3 0 1 0 -1E6
E24 4 0 2 0 -1E6

G14 1 4 0 31 32.000M
R14 31 0 1000
T14 30 0 31 0 Z0=1000 TD=1.0000U
E14 30 0 1 4 1

G23 2 3 0 41 32.000M
R23 41 0 1000
T23 40 0 41 0 Z0=1000 TD=1.0000U
E23 40 0 2 3 1

.ENDS
.AC DEC 50 1K 500K
.OPTIONS PIVTOL=1E-20 LIMPTS=20000
*.TRAN .05U 50U
 
*ALIAS  V(12)=VOUT
.PRINT AC  V(12)  VP(12)  V(4)  VP(4) 
.PRINT TRAN  V(12) 
X4 12 2 CRES#0  
*{C=2P } 
X5 39 2 CRES#0  
*{C=2P } 
X8 4 6 NSTR#0  
*{TD=1U C=2P } 
X9 3 6 12 9 ZINT#0  
*{TD=1U C=32P } 
E1 11 0 0 10 20K
R1 10 4 100K
R2 10 11 10K
V1 39 0 PULSE 0 2 AC 1
X11 11 2 NSTR#0  
*{TD=1U C=2P } 
X2 2 5 4 8 ZINT#0  
*{TD=1U C=32P } 
.END