scn5
*SPICE_NET
.AC DEC 50 1K 500K
.OPTIONS ACCT PIVTOL=1E-20 LIMPTS=10000
.TRAN 1U 20U 
*INCLUDE SCN.LIB
.SUBCKT ZINT#0 1 2 3 4 
* 2 PHASE INT, 1 3 ARE ODD IN->OUT; 2,4 ARE EVEN
R1 1 3 31.250 
R2 2 4 31.250 
E13 3 0 1 0 -1E6
E24 4 0 2 0 -1E6
G14 1 4 0 31 32.000M
R14 31 0 1000
T14 30 0 31 0 Z0=1000 TD=1.0000U
E14 30 0 1 4 1
G23 2 3 0 41 32.000M
R23 41 0 1000
T23 40 0 41 0 Z0=1000 TD=1.0000U
E23 40 0 2 3 1
.ENDS
.SUBCKT CRES#0 1 2
R1 1 2 500.00 
.ENDS
.SUBCKT NSTR#0 1 2
*NEGATIVE STORISTER I = 1E9 * (- C * Z^-1/2)
E1 3 0 1 2 1
T1 3 0 4 0 Z0=1000 TD=1.0000U
RT 4 0 1000
G1 1 2 0 4 2.0000M
.ENDS
.SUBCKT SCNAMP  2    3  6   
*             - IN   +  OUT 
*DERIVED FROM OPAMP IN LIN.LIB
*
RIP 3 0 10MEG
CIP 3 0 1.4PF
IBN 2 0 1.0000P
RIN 2 0 10MEG
CIN 2 0 1.4PF
VOFST 2 10 
RID 10 3 200K
EA 11 0 10 3 1
R1 11 12 5K
R2 12 13 50K
C1 12 0 5.2000P
GA 0 14 0 13 378.00 
C2 13 14 1.0800P
RO 14 0 75
L 14 6 12.000U
RL 14 6 1000
CL 6 0 3PF
.ENDS
.SUBCKT MF10HZ100 15  4    3   2   5   20  19  16  1   18  17 
*Connections   AGND INVA HPA BPA S1A LPB BPB S1B LPA HPB INVB
*FOR GAIN OF 100 DEFINE 2P=2P, 
*FOR GAIN OF 50 DEFINE 2P=4P
*DEFINE /SCNCAP=2P
X19 31 30 19 34 ZINT#0  
*{TD=1U C=32P } 
X2 35 36 2 33 ZINT#0  
*{TD=1U C=32P } 
X4 1 35 CRES#0  
*{C= 2P } 
X5 5 35 CRES#0  
*{C= 2P } 
X8 2 29 NSTR#0  
*{TD=1U C= 2P } 
X9 28 29 1 32 ZINT#0  
*{TD=1U C=32P } 
XE1 4 15 3 SCNAMP
X11 3 35 NSTR#0  
*{TD=1U C= 2P } 
X20 20 31 CRES#0  
*{C= 2P } 
X21 16 31 CRES#0  
*{C= 2P } 
X22 19 38 NSTR#0  
*{TD=1U C= 2P } 
X23 37 38 20 40 ZINT#0  
*{TD=1U C=32P } 
X24 18 31 NSTR#0  
*{TD=1U C= 2P } 
XE2 17 15 18 SCNAMP
.ENDS
*INCLUDE SYS.LIB
*ALIAS  V(4)=VOUTA
*ALIAS  V(2)=VOUTB
.PRINT AC  V(4)  VP(4)  V(2)  VP(2) 
.PRINT TRAN  V(4)  V(2) 
R2 11 12 100K
R3 14 15 10K
R4 14 16 100K
V1 3 0 PULSE 0 2 AC 1
V2 1 0 PULSE 0 2 AC 1
X9 0 11 10 12 1 2 16 3 4 15 14 MF10HZ10 
R1 11 10 10K
.END