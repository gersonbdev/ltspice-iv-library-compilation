scn6
*SPICE_NET
*INCLUDE SYS.LIB
*INCLUDE SCN.LIB
X12 6 11 13 MUL  {K=1 } 
X13 19 11 22 MUL  {K=1 } 
X15 13 19 SINT  {K=31.25K } 
X16 22 20 SINT  {K=31.25K } 
X17 3 3 1 SCNAMP2 
X18 20 4 16 7 SUM3  {K1=-1 K2=1 K3=-1 } 
X19 7 8 9 MUL  {K=1 } 
X20 19 8 14 MUL  {K=1 } 
X21 9 19 SINT  {K=31.25K } 
X22 14 20 SINT  {K=31.25K } 
X23 10 12 4 SCNAMP2 
X14 3 1 16 6 SUM3  {K1=-1 K2=1 K3=-1 } 
.END