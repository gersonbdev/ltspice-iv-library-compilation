IBIS
*SPICE_NET
.TRAN .1N 120N
*INCLUDE IBIS1.LIB
.OPTION ACCT VSCALE=7.5
*ALIAS  V(100)=VINPUT
*ALIAS  V(500)=ENABLE
*ALIAS  V(1)=VB
*ALIAS  V(14)=VA
*ALIAS  V(3)=VLOAD2
*ALIAS  V(17)=VLOAD10
.PRINT TRAN  V(100)  V(500)  V(1)  V(14) 
.PRINT TRAN  V(3)  V(17) 
X36 3 300 400 PCIIW
V1 100 0 PULSE 0 5 0 2.5N 2.5N 30N 60N
V2 500 0 5
V3 300 0 5.25
V4 400 0 0
X6 100 14 300 400 500 PCIOW
X16 100 1 300 400 500 PCIOW
C1 1 0 40PF
X32 9 300 400 PCIIW
X33 22 300 400 PCIIW
X34 23 300 400 PCIIW
X35 24 300 400 PCIIW
X37 6 300 400 PCIIW
X38 4 300 400 PCIIW
X39 8 300 400 PCIIW
C2 11 0 .5PF
C3 10 0 .5PF
C4 5 0 .5PF
C5 16 0 .5PF
C6 15 0 .5PF
C7 7 0 .5PF
C8 13 0 .5PF
C9 12 0 .5PF
C10 18 0 .5PF
X3 14 11 BLINE {LENGTH=1 }
X97 11 7 BLINE {LENGTH=1 }
X98 7 10 BLINE {LENGTH=1 }
X99 10 13 BLINE {LENGTH=1 }
X100 13 5 BLINE {LENGTH=1 }
X101 5 12 BLINE {LENGTH=1 }
X102 12 16 BLINE {LENGTH=1 }
X103 16 18 BLINE {LENGTH=1 }
X104 18 15 BLINE {LENGTH=1 }
X105 3 11 BLINE1 {LENGTH=1.5 }
X106 6 10 BLINE1 {LENGTH=1.5 }
X107 4 5 BLINE1 {LENGTH=1.5 }
X108 8 16 BLINE1 {LENGTH=1.5 }
X109 17 15 BLINE1 {LENGTH=1.5 }
X110 9 7 BLINE1 {LENGTH=1.5 }
X111 22 13 BLINE1 {LENGTH=1.5 }
X112 23 12 BLINE1 {LENGTH=1.5 }
X113 24 18 BLINE1 {LENGTH=1.5 }
X40 17 300 400 PCIIW
.END
