IBIS
*SPICE_NET
*dEFINE RTF=34K
*dEFINE RTR=31K
.TRAN .1N 50N
*INCLUDE INTEL.LIB
.SUBCKT EPWL_DN  3    4    1   2
*               out+ OUT- IN+ IN-
	B1 3 4 V= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + -109.99999M :
+ (V(1,2) < -4.0000000) ? 2.9999999M*V(1,2) + -94.999995M :
+ (V(1,2) < -3.0000000) ? 3.9999998M*V(1,2) + -90.999996M :
+ (V(1,2) < -2.0000000) ? 11.999999M*V(1,2) + -66.999997M :
+ (V(1,2) < -1.0000000) ? 33.999998M*V(1,2) + -22.999999M :
+ (V(1,2) < 0.0000000E+00) ? 56.999997M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 499.99998M) ? 61.999997M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 1.0000000) ? 51.999998M*V(1,2) + 4.9999998M :
+ (V(1,2) < 1.5000000) ? 37.999998M*V(1,2) + 18.999999M :
+ (V(1,2) < 2.0000000) ? 29.999999M*V(1,2) + 30.999999M :
+ (V(1,2) < 2.5000000) ? 17.999999M*V(1,2) + 54.999997M :
+ (V(1,2) < 3.0000000) ? 5.9999997M*V(1,2) + 84.999996M :
+ (V(1,2) < 3.5000000) ? 3.9999998M*V(1,2) + 90.999996M :
+ (V(1,2) < 4.0000000) ? 3.9999998M*V(1,2) + 90.999996M :
+ (V(1,2) < 4.5000000) ? 3.9999998M*V(1,2) + 90.999996M :
+ (V(1,2) < 5.0000000) ? 3.9999998M*V(1,2) + 90.999996M :
+ (V(1,2) < 10.0000000) ? 1.7999999M*V(1,2) + 102.00000M :
+ 1.0000000N*V(1,2) + 119.99998M
.ENDS
.SUBCKT EPWL_UP 3    4    1   2
*               out+ OUT- IN+ IN-
	B1 3 4 V= 
+ (V(1,2) < -5.0000000) ? -1.0000000N*V(1,2) + 56.999992M :
+ (V(1,2) < -4.0000000) ? -2.9999999M*V(1,2) + 41.999998M :
+ (V(1,2) < -3.0000000) ? -3.9999998M*V(1,2) + 37.999998M :
+ (V(1,2) < -2.0000000) ? -9.9999995M*V(1,2) + 19.999999M :
+ (V(1,2) < -1.0000000) ? -16.999999M*V(1,2) + 5.9999997M :
+ (V(1,2) < 0.0000000E+00) ? -22.999999M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 499.99998M) ? -25.999999M*V(1,2) + 0.0000000E+00 :
+ (V(1,2) < 1.0000000) ? -19.999999M*V(1,2) + -2.9999999M :
+ (V(1,2) < 1.5000000) ? -19.999999M*V(1,2) + -2.9999999M :
+ (V(1,2) < 2.0000000) ? -13.999999M*V(1,2) + -11.999999M :
+ (V(1,2) < 2.5000000) ? -11.999999M*V(1,2) + -15.999999M :
+ (V(1,2) < 3.0000000) ? -7.9999996M*V(1,2) + -25.999999M :
+ (V(1,2) < 3.5000000) ? -3.9999998M*V(1,2) + -37.999998M :
+ (V(1,2) < 4.5000000) ? -2.9999999M*V(1,2) + -41.499998M :
+ (V(1,2) < 5.0000000) ? -3.9999998M*V(1,2) + -36.999998M :
+ (V(1,2) < 10.0000000) ? -1.7999999M*V(1,2) + -47.999998M :
+ -1.0000000N*V(1,2) + -65.999987M
.ENDS
.SUBCKT VCC_OUT 3    4    1   2
*               out+ OUT- IN+ IN-
B1 3 4 I= 
+ (V(1,2) < 5.6000000) ? -1.0000000N*V(1,2) + 5.6000002N :
+ (V(1,2) < 5.7000000) ? 39.999998M*V(1,2) + -223.99999M :
+ (V(1,2) < 5.8000000) ? 259.99999M*V(1,2) + -1.4780000 :
+ (V(1,2) < 5.9000000) ? 219.99999M*V(1,2) + -1.2460000 :
+ (V(1,2) < 6.0000000) ? 219.99999M*V(1,2) + -1.2460000 :
+ (V(1,2) < 10.0000000) ? 223.99999M*V(1,2) + -1.2700000 :
+ -1.0000000N*V(1,2) + 969.99996M
.ENDS
.SUBCKT GND_OUT  3    4    1   2
*               out+ OUT- IN+ IN-
B1 3 4 I= 
+ (V(1,2) < -5.0000000) ? 1.0000000N*V(1,2) + -1.7250000 :
+ (V(1,2) < -1.0000000) ? 403.74998M*V(1,2) + 293.74999M :
+ (V(1,2) < -899.99996M) ? 399.99998M*V(1,2) + 289.99999M :
+ (V(1,2) < -799.99996M) ? 349.99998M*V(1,2) + 244.99999M :
+ (V(1,2) < -699.99997M) ? 299.99999M*V(1,2) + 204.99999M :
+ (V(1,2) < -599.99997M) ? 49.999998M*V(1,2) + 29.999999M :
+ 1.0000000N*V(1,2) + 600.00000P
.ENDS
.OPTIONS ACCT 
*ALIAS  V(220)=VOUT
*ALIAS  V(850)=VRUP
*ALIAS  V(4)=VOUT
*ALIAS  I(V5)=IDIE
*ALIAS  I(V6)=IINT2
*ALIAS  I(V7)=IINT1
.PRINT TRAN  V(220)  V(840)  V(850)  V(100) 
.PRINT TRAN  V(500)  V(830)  V(820)  V(4) 
.PRINT TRAN  I(V5) I(V6) I(V7)
B1 820 0 V=V(100) & V(500)
B2 830 0 V= V(500) & ~V(100)
S1 220 850 0 820 SMOD
.MODEL SMOD SW RON=.1M ROFF=1E15 VT=-1.2 VH=.1
S2 840 220 0 830 SMOD
C1 300 850 .01P
C2 840 400 .01P
V1 100 0 PULSE 0 5 0 0 0 10N 20N
V2 500 0 PULSE 0 5 0 0 0 5N 10N
V3 300 0 5
V4 400 0 0
B3 300 850 I= V(830) > 1.2   ? 0 : V(300,850) / 31K
B4 840 400 I= V(820) > 1.2 ? 0 : V(840,400) / 34K
XEPL_DN 2 400 8 840 EPWL_DN
G1 8 400 2 8 1
R1 6 400 1
X1 3 300 850 8 EPWL_UP
G2 300 8 8 3 1
R2 300 6 1
XVCC_OUT 6 300 300 6 VCC_OUT
XGND_OUT 6 400 6 400 GND_OUT
R3 5 1 100
R4 1 4 .277
C3 4 400 1.36P
C4 5 400 5.64P
L1 5 1 32.75N
V5 6 5 
V6 8 6 
V7 220 8 
.END
