SCN14
.OPTIONS LIMPTS=1000
*SPICE_NET
*INCLUDE SCN.LIB
.SUBCKT SCNAMP64 2    3  6
*                - IN + OUT
*PARAMS ARE GAIN=80.000  FT=7.0000MEG IOS=1.0000P VOS=1.0000M IBIAS=3.0000P     
*GAIN IS IN db  
RIP 3 0 10MEG   
CIP 3 0 1.4PF   
IBN 2 0 3.0000P 
RIN 2 0 10MEG   
CIN 2 0 1.4PF   
VOFST 2 10 1.0000M      
RID 10 3 200K   
EA 11 0 10 3 1  
R1 11 12 5K     
R2 12 13 50K    
C1 12 0 1.8571P 
GA 0 14 0 13 135.00     
C2 13 14 385.71F
RO 14 0 75      
L 14 6 4.2857U  
RL 14 6 1000    
CL 6 0 3PF      
.ENDS   
.SUBCKT LT6410D 3 2 1 33 28 10 4 6 14 29 12 5 22 24 30 13 8 31 32 26 17
*Connections   INVA AGND HPA SA BPA LPA INVB HPB SB BPB LPB 
*Connections                    INVC HPC SC BPC LPC INVD HPD BPD LPD CLK
* Subcircuit for DIP package
X10 16 17 18 MUL#0  
*{K=1 } 
X11 28 17 20 MUL#0  
*{K=1 } 
X12 18 28 SINT#0  
*{K=31.25K } 
X13 20 10 SINT#0  
*{K=31.25K } 
X15 1 33 16 SUM2#0  
*{K1=1 K2=-1 }
X16 4 2 6 SCNAMP64
X17 7 17 9 MUL#0  
*{K=1 } 
X18 29 17 11 MUL#0  
*{K=1 } 
X19 9 29 SINT#0  
*{K=31.25K } 
X20 11 12 SINT#0  
*{K=31.25K } 
X21 6 14 7 SUM2#0  
*{K1=1 K2=-1 }
X22 5 2 22 SCNAMP64
X23 23 17 25 MUL#0  
*{K=1 } 
X24 30 17 27 MUL#0  
*{K=1 } 
X25 25 30 SINT#0  
*{K=31.25K } 
X26 27 13 SINT#0  
*{K=31.25K } 
X27 22 24 23 SUM2#0  
*{K1=1 K2=-1 }
X28 8 2 31 SCNAMP64
X29 31 17 34 MUL#0  
*{K=1 } 
X30 32 17 36 MUL#0  
*{K=1 } 
X31 34 32 SINT#0  
*{K=31.25K } 
X32 36 26 SINT#0  
*{K=31.25K } 
X5 3 2 1 SCNAMP64
.ENDS
*INCLUDE SYS.LIB
.SUBCKT MUL#0 1 2 3
RIN1 1 0 1E12
RIN2 2 0 1E12
ROUT 3 0 1E12
E1 3 0 POLY(2) 1 0 2 0 0 0 0 0 1.0000 
.ENDS
.SUBCKT SINT#0 1 2
*PARAMS ARE GAIN=31.250K
RIN 1 0 1E12
E1 3 0 0 1 31.250K
C1 2 4 1U IC=0
R1 3 4 1MEG
E2 2 0 0 4 1.0000MEG
.ENDS
.SUBCKT SUM2#0 1 2 3
RIN1 1 0 1E12
RIN2 2 0 1E12
ROUT 3 0 1E12
E1 3 0 POLY(2) 1 0 2 0 0 1.0000  -1.0000 
.ENDS
.AC DEC 10 1K 10MEG
*ALIAS  V(19)=VOUT
.PRINT AC  V(19)  VP(19) 
R73 2 3 100.86K
R74 19 5 25.42K
R75 6 5 17.72K
R76 7 5 11.52K
V14 3 0 AC 1
R77 8 9 99.83K
R78 10 9 68.15K
R79 11 9 10.18K
R80 8 5 13.84K
R82 12 9 16.61K
R84 13 14 20.93K
R85 15 14 45.2K
R86 12 14 25.52K
R87 14 16 25.72K
R88 2 17 99.73K
R89 2 16 23.6K
R90 2 18 16.75K
X8 2 0 18 0 16 17 14 13 0 15 12 9 11 8 10 8 5 7 6 19 1 LT6410D 
V13 1 0 10
.END