*** SAMTEC MODEL TEST FILE 
** 2 rows 10 pins each row x 8 section
** for 50 ps edge rate or slower
*     
* column*01*02*03*04*05*06*07*08*09*10
* row A...X  X  X  A  X  X  X  X  X  X
* ground..X 
* row B...X  X  X  X  X  X  X  X  X  X
* "X=REF, A=ACTIVE"     
* "Q=QUIET, M=MONITORED"     
*     
*************************************     
*     
* QTS-RA QSS-01
* 1.0V/50PS TR  
* 50 OHM TERMINATIONS  
*   
*   
******* input/output instructions *************  
* driven lines  
.PRINT TRAN V(1104) V(3104)
* quiet lines  
.PRINT TRAN V(1103) V(3103)
********** analysis & control ***************** 
.OPTIONS METHOD=GEAR RELTOL=.001
.TRAN 5PS 1NS  
************** excitation *********************  
XDR1 1104 0 SRC50PS  
XDR2 1304 0 SRC50PS
*   
************** analysis & control *************** 
********************************   
.SUBCKT SRC50PS 3 2
*1.0v; 50ps; 20-80% 
********************  
VS1 1 2 PWL(
+0 0
+.02NS 0.06 
+.03NS 0.14 
+.04NS 0.24 
+.05NS 0.4 
+.1NS 1.6 
+.11NS 1.76 
+.12NS 1.86 
+.13NS 1.94 
+.15NS 2) 
RS1 1 3 50
************  
.ENDS SRC50PS 
************  
********************************  
.SUBCKT SRC100PS 3 2
*1.0v; 100ps; 20-80% 
********************  
VS1 1 2 PWL(
+0 0
+.04NS 0.06 
+.06NS 0.14 
+.08NS 0.24 
+.1NS 0.4 
+.2NS 1.6 
+.22NS 1.76 
+.24NS 1.86 
+.26NS 1.94 
+.3NS 2) 
RS1 1 3 50
************  
.ENDS SRC100PS 
************  
********************************  
.SUBCKT SRC500PS 3 2
*1.0v; 0.5NS; 20-80% 
********************  
VS1 1 2 PWL(
+0 0
+.2NS 0.06 
+.3NS 0.14 
+.4NS 0.24 
+.5NS 0.4 
+1NS 1.6 
+1.1NS 1.76 
+1.2NS 1.86 
+1.3NS 1.94 
+1.5NS 2) 
RS1 1 3 50
************  
.ENDS SRC500PS 
********************************  
.SUBCKT SRC1000PS 3 2
*1.0v; 1NS; 20-80% 
********************  
VS1 1 2 PWL(
+0 0
+.4NS 0.06 
+.6NS 0.14 
+.8NS 0.24 
+1NS 0.4 
+2NS 1.6 
+2.2NS 1.76 
+2.4NS 1.86 
+2.6NS 1.94 
+3NS 2) 
RS1 1 3 50
************  
.ENDS SRC1000PS 
************  
.SUBCKT ACDR11 1 3
V1 1 2 AC
R1 2 3 50
.ENDS ACDR11
********************************END OF DRIVERS 
**side a********** 
*  
RR1101 1101 0 .001
RR1102 1102 0 .001
RR1103 1103 0 .001
*RR1104 1104 0 .001
RR1105 1105 0 .001
RR1106 1106 0 .001
RR1107 1107 0 .001
RR1108 1108 0 .001
RR1109 1109 0 .001
RR1110 1110 0 .001
*
************** reference ********************* 
RR1201 1201 0 .001
*  
**side b********** 
RR1301 1301 0 .001
RR1302 1302 0 .001
RR1303 1303 0 .001
*RR1304 1304 0 .001
RR1305 1305 0 .001
RR1306 1306 0 .001
RR1307 1307 0 .001
RR1308 1308 0 .001
RR1309 1309 0 .001
RR1310 1310 0 .001
*  
**side a********** 
*  
RR3101 3101 0 .001
RR3102 3102 0 .001
RR3103 3103 0 .001
*RR3104 3104 0 .001
RR3105 3105 0 .001
RR3106 3106 0 .001
RR3107 3107 0 .001
RR3108 3108 0 .001
RR3109 3109 0 .001
RR3110 3110 0 .001
*
************** referencing ******************** 
RR3201 3201 0 .001
*  
**side b********** 
RR3301 3301 0 .001
RR3302 3302 0 .001
RR3303 3303 0 .001
*RR3304 3304 0 .001
RR3305 3305 0 .001
RR3306 3306 0 .001
RR3307 3307 0 .001
RR3308 3308 0 .001
RR3309 3309 0 .001
RR3310 3310 0 .001
*  
************* terminations ******************** 
*  
** side a ******
*  
RT1101 1101 0 50
RT1102 1102 0 50
RT1103 1103 0 50
*RT1104 1104 0 50
RT1105 1105 0 50
RT1106 1106 0 50
RT1107 1107 0 50
RT1108 1108 0 50
RT1109 1109 0 50
RT1110 1110 0 50
*  
**side b********** 
*  
RT1301 1301 0 50
RT1302 1302 0 50
RT1303 1303 0 50
*RT1304 1304 0 50
RT1305 1305 0 50
RT1306 1306 0 50
RT1307 1307 0 50
RT1308 1308 0 50
RT1309 1309 0 50
RT1310 1310 0 50
*  
** side a ******
*  
RT3101 3101 0 50
RT3102 3102 0 50
RT3103 3103 0 50
RT3104 3104 0 50
RT3105 3105 0 50
RT3106 3106 0 50
RT3107 3107 0 50
RT3108 3108 0 50
RT3109 3109 0 50
RT3110 3110 0 50
*  
**side b********** 
*  
RT3301 3301 0 50
RT3302 3302 0 50
RT3303 3303 0 50
RT3304 3304 0 50
RT3305 3305 0 50
RT3306 3306 0 50
RT3307 3307 0 50
RT3308 3308 0 50
RT3309 3309 0 50
RT3310 3310 0 50
*  
* PCB PAD CAPACITANCE
** side a *********
*  
CP1101 1101 0 .1PF
CP1102 1102 0 .1PF
CP1103 1103 0 .1PF
CP1104 1104 0 .1PF
CP1105 1105 0 .1PF
CP1106 1106 0 .1PF
CP1107 1107 0 .1PF
CP1108 1108 0 .1PF
CP1109 1109 0 .1PF
CP1110 1110 0 .1PF
*  
** side b ******
*  
CP1301 1301 0 .1PF
CP1302 1302 0 .1PF
CP1303 1303 0 .1PF
CP1304 1304 0 .1PF
CP1305 1305 0 .1PF
CP1306 1306 0 .1PF
CP1307 1307 0 .1PF
CP1308 1308 0 .1PF
CP1309 1309 0 .1PF
CP1310 1310 0 .1PF
*  
** side a *********
*  
CP3101 3101 0 .1PF
CP3102 3102 0 .1PF
CP3103 3103 0 .1PF
CP3104 3104 0 .1PF
CP3105 3105 0 .1PF
CP3106 3106 0 .1PF
CP3107 3107 0 .1PF
CP3108 3108 0 .1PF
CP3109 3109 0 .1PF
CP3110 3110 0 .1PF
*  
** side b ******
*  
CP3301 3301 0 .1PF
CP3302 3302 0 .1PF
CP3303 3303 0 .1PF
CP3304 3304 0 .1PF
CP3305 3305 0 .1PF
CP3306 3306 0 .1PF
CP3307 3307 0 .1PF
CP3308 3308 0 .1PF
CP3309 3309 0 .1PF
CP3310 3310 0 .1PF
*  
*  
*******************   
*   
XC
* outer
+ 1101 1102 1103 1104 1105 1106 1107 1108
* ground ******************************************
+ 1201
* inner
+ 1301 1302 1303 1304 1305 1306 1307 1308
* BEVEL * QSS *************************************
* outer row ***************************************
+ 3101 3102 3103 3104 3105 3106 3107 3108
* ground ******************************************
+ 3201
* inner row ***************************************
+ 3301 3302 3303 3304 3305 3306 3307 3308
+ QTSRAQSS
********
.INCLUDE m_qtsra_qss01.cir
********   
.END
