*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Inc.
* Models developed and under copyright by:
* National Semiconductor, Inc.  

*/////////////////////////////////////////////////////////////////////
* Legal Notice: This material is intended for free software support.
* The file may be copied, and distributed; however, reselling the 
*  material is illegal

*////////////////////////////////////////////////////////////////////
* For ordering or technical information on these models, contact:
* National Semiconductor's Customer Response Center
*                 7:00 A.M.--7:00 P.M.  U.S. Central Time
*                                (800) 272-9959
* For Applications support, contact the Internet address:
*  amps-apps@galaxy.nsc.com

*//////////////////////////////////////////////////////////
*LM6118 Fast Settling Dual OP-AMP MACRO-MODEL
*//////////////////////////////////////////////////////////
*
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   positive power supply
*                   |   |   |   negative power supply
*                   |   |   |   |   output
*                   |   |   |   |   |
*                   |   |   |   |   |
.SUBCKT LM6118/NS   1   2  99  50  28
*
*Features:
*Low offset voltage =   .2mV
*High bandwidth =      17MHz
*Slew rate (Av=-1) = 140V/uS
*
*NOTE: Model is for single device only and simulated
*      supply current is 1/2 of total device current.
*
****************INPUT STAGE**************
*
IOS 2 1 20N
*^Input offset current
CI1 1 0 2.5P
CI2 2 0 2.5P
R1  1 3 3.125G
R2  3 2 3.125G
I1 99 4 40U
R43 45 4 1.25K
R44 46 4 1.25K
Q1  5 2 45 QX
Q2  6 7 46 QX
R3 50 5 2.54K
R4 50 6 2.54K
*Fp2=30 MHz
C4 5 6 1.0433P
*
***********COMMON MODE EFFECT***********
*
I2 99 50 2.71M
*^Quiescent supply current
EOS 7 1 POLY(1) 16 49 .2E-3 1
*Input offset voltage.^
R8 99 49 71.4K
R9 49 50 71.4K
*
*********OUTPUT VOLTAGE LIMITING********
V2 99 8 2.63
D1 9 8 DX
D2 10 9 DX
V3 10 50 2.63
*
**************SECOND STAGE**************
*
EH 99 98 99 49 1
G1 98 9 POLY(1) 5 6 0 5E-3 0 5.056
*Fp1=38.24 Hz
R5 98 9 100MEG
C3 98 9 41.62P
*
***************POLE STAGE***************
*
*Fp=110 MHz
G3 98 15 9 49 1E-6
R12 98 15 1MEG
C5 98 15 1.4469E-15
*
*********COMMON-MODE ZERO STAGE*********
*
*Fpcm=6 KHz
G4 98 16 3 49 1E-8
L2 98 17 26.526M
R13 17 16 1K
*
**************OUTPUT STAGE**************
*
F6 50 99 POLY(1) V6 200U 1
E1 99 23 99 15 1
R16 24 23 10
D5 26 24 DY
V6 26 22 .63V
R17 23 25 10
D6 25 27 DY
C9 23 22 .001U
V7 22 27 .63V
V5 22 21 .63V
D4 21 15 DX
V4 20 22 .63V
D3 15 20 DX
L3 22 28 100P
RL3 22 28 100K
*
***************MODELS USED**************
*
.MODEL DX D(IS=1E-15)
.MODEL DY D(IS=1E-25)
.MODEL QX PNP(BF=100)
*
.ENDS
*$
