scn5
*SPICE_NET
.AC DEC 50 1K 500K
.OPTIONS ACCT PIVTOL=1E-20 LIMPTS=10000
.TRAN 1U 20U 
*INCLUDE SCN.LIB
*ALIAS  V(4)=VOUTA
*ALIAS  V(2)=VOUTB
.PRINT AC  V(4)  VP(4)  V(2)  VP(2) 
.PRINT TRAN  V(4)  V(2) 
R2 11 12 100K
R3 14 15 10K
R4 14 16 100K
V1 3 0 PULSE 0 2 AC 1
V2 1 0 PULSE 0 2 AC 1
X9 0 11 10 12 1 2 16 3 4 15 14 MF10HZ10 
R1 11 10 10K
.END