IBIS
*SPICE_NET
.TRAN .1N 120N
*INCLUDE IBIS1.LIB
.OPTION ACCT VSCALE=5
*INCLUDE FRAME.LIB
*ALIAS  V(100)=VINPUT
*ALIAS  V(500)=ENABLE
*ALIAS  V(7)=VOUT
.PRINT TRAN  V(100)  V(500)  V(7) 
V2 500 0 5
V3 300 0 5
V4 400 0 0
X6 100 7 300 400 500 PCIOW
C1 7 0 50PF
V1 100 0 PULSE 0 5 0 2.5N 2.5N 27.44N 59.88N
.END
