IBIS
*SPICE_NET
*DEFINE RTF=34K
*DEFINE RTR=31K
.TRAN .1N 50N
*INCLUDE INTEL.LIB
.OPTIONS ACCT 
*ALIAS  V(220)=VOUT
*ALIAS  V(850)=VRUP
*ALIAS  V(4)=VOUT
*ALIAS  I(V5)=IDIE
*ALIAS  I(V6)=IINT2
*ALIAS  I(V7)=IINT1
.PRINT TRAN  V(220)  V(840)  V(850)  V(100) 
.PRINT TRAN  V(500)  V(830)  V(820)  V(4) 
.PRINT TRAN  I(V5) I(V6) I(V7)
B1 820 0 V=V(100) & V(500)
B2 830 0 V= V(500) & ~V(100)
S1 220 850 0 820 SMOD
.MODEL SMOD SW RON=.1M ROFF=1E15 VT=-1.2 VH=.1
S2 840 220 0 830 SMOD
C1 300 850 .01P
C2 840 400 .01P
V1 100 0 PULSE 0 5 0 0 0 10N 20N
V2 500 0 PULSE 0 5 0 0 0 5N 10N
V3 300 0 5
V4 400 0 0
B3 300 850 I= V(830) > 1.2   ? 0 : V(300,850) / RTR
B4 840 400 I= V(820) > 1.2 ? 0 : V(840,400) / RTF
XEPL_DN 2 400 8 840 EPWL_DN
G1 8 400 2 8 1
R1 6 400 1
X1 3 300 850 8 EPWL_UP
G2 300 8 8 3 1
R2 300 6 1
XVCC_OUT 6 300 300 6 VCC_OUT
XGND_OUT 6 400 6 400 GND_OUT
R3 5 1 100
R4 1 4 .277
C3 4 400 1.36P
C4 5 400 5.64P
L1 5 1 32.75N
V5 6 5 
V6 8 6 
V7 220 8 
.END
