555_TIMER1.CIR - ASTABLE MODE
*
VCC	1	0	5V
*
* EXTERNAL TIMING COMPONENTS
RA	1	2	1K
RB	2	3	10K
C1	3	0	100PF
*
* DISCHARGE TRANSISTOR
Q1	2 6 0	QNOM
RBQ	15	6	15K
*
* 1/3 AND 2/3 VCC DIVIDER
R1	1	4	5K
R2	4	5	5K
R3	5	0	5K
*
* COMPARATORS
XCMP1	3 4 11 COMP1 
XCMP2	5 3 12 COMP1 
*
* RS FLIP-FLOP
XNOT1	11 13 1 NOT
XNOT2	12 16 1 NOT
XNAND1	13 14 15 1	NAND
XNAND2	15 16 14 1	NAND
*
* SUBCIRCUITS AND MODELS ***********************************
*
.SUBCKT NAND 1 2 3 4
* TERMINALS A B OUT VCC
RL	3	4	500
CL	3	0	10PF
S1	3 5	1 0 	SW
S2	5 0	2 0 	SW
.ENDS
*
.SUBCKT NOT 1 3 4
* TERMINALS A OUT VCC
RL	3	4	500
CL	3	0	10PF
S1	3 0	1 0 	SW
.ENDS
*
*
.SUBCKT COMP1  1 2 5
* TERMINALS: 1-INPUT+, 2-INPUT-, 5-OUTPUT
* DIFF AMP WITH HYSTERESIS
EDIFF	3	0	VALUE = { V(1) - V(2) + V(5)/500 }
* FREQUENCY RESPONSE
RP1	3	4	200
CP1	4	0	100PF
* LIMITER
EOUT	5	0	TABLE {V(4)} = (-1MV 0V) (1MV, 5V) 
.ENDS
*
*
.MODEL	SW	VSWITCH(VON=3 VOFF=2 RON=10 ROFF=100K)
.model	QNOM	NPN(BF=100)
*
* ANALYSIS *************************************************
.TRAN 	0.05US  5US UIC
.IC V(15)=0V V(14)=5V V(3)=0V
*
* VIEW RESULTS *********************************************
.PRINT	TRAN 	V(3) V(14)
.PROBE
.END