*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Inc.
* Models developed and under copyright by:
* National Semiconductor, Inc.  

*/////////////////////////////////////////////////////////////////////
* Legal Notice: This material is intended for free software support.
* The file may be copied, and distributed; however, reselling the 
*  material is illegal

*////////////////////////////////////////////////////////////////////
* For ordering or technical information on these models, contact:
* National Semiconductor's Customer Response Center
*                 7:00 A.M.--7:00 P.M.  U.S. Central Time
*                                (800) 272-9959
* For Applications support, contact the Internet address:
*  Appshelp@galaxy.nsc.com

*/////////////////////////////////////////////////
*LM6311 Operational Amplifier Macro-Model
*/////////////////////////////////////////////////
*
* Connections:     Non-Inverting Input
*                  | Inverting
*                  | | Output
*                  | | | +Vcc
*                  | | | | -Vee
*                  | | | | | External Compensation
*                  | | | | | | 
*                  | | | | | | 
.SUBCKT LM6311/NS 3 2 6 7 4 5 
*Features
*   This is an Ultra Low Noise, Wideband Monolithic Voltage
*   Feedback Op Amp with Current Supply Adjust and External
*   Compensation.
*
*
* BIAS CIRCUITRY
*
R1 7 10 100
Q1 10 12 11 QINN1
D1 11 12 DZ
R2 11 8 1.00K
C1 8 0 1.00P
R3 8 4 1.00G
R4 7 12 100K
D2 12 13 DZ
D3 13 4 DZ
*
G1 0 14 POLY(3) 12 4  7 10 0 14 -226M 294M -10.0 1.00M
D4 0 14 DY
*
G2 7 20 POLY(2) 14 0 7 20 -442N 2.56U 1.39U
C2 20 0 800F
G7 7 34 POLY(2) 14 0 7 34 -442N 2.56U 1.39U
C5 34 0 800F
*
G4 21 4 POLY(2) 14 0 21 4 9.27U 5.43U 400N
C4 21 0 400F
G9 36 4 POLY(2) 14 0 36 4 9.27U 5.43U 400N
C7 36 0 400F
*
* INPUT STAGE
*
C3 2 0 1.00P
G3 2 0 POLY(2) 50 0 51 0 0 100U 100U
Q2 4 2 20 QINP2
Q3 7 2 21 QINN1
V1 7 22 DC 1.00
Q4 22 20 23 QINN1
Q5 24 21 23 QINP2
V2 24 4 DC 1.00
*
Q6 31 34 23 QINN2
Q7 32 36 23 QINP1
Q8 7 35 36 QINN2
Q9 4 35 34 QINP1
G8 35 0 POLY(2) 52 0 53 0 0 100U 100U
E1 3 35 POLY(2) 54 0 55 0 1.55M 1.00 1.00
C6 3 0 1.00P
*
* GAIN STAGE
*
D5 7 30 DY
G5 30 31 POLY(1) 30 31 0 1.00
R5 7 31 450
V3 7 40 DC 1.75
D7 41 40 DX
C8 7 41 7.00P
G10 7 41 POLY(3) 7 41 7 31 30 31 0 574N 2.22M 250M 0 4.78U 538U
C11 31 43 400F
G12 7 43 POLY(1) 7 31 0 2.22M
C12 43 0 800F
*
G6 32 33 POLY(1) 32 33 0 1.00
D6 33 4 DY
R6 32 4 450
D8 42 41 DX
V4 42 4 DC 1.75
C10 41 4 7.00P
G11 41 4 POLY(3) 41 4 32 4 32 33 0 1.33U 2.22M 250M 0 11.1U 1.25M
C13 32 44 800F
G13 44 4 POLY(1) 32 4 0 8.00M
C14 44 0 400F
*
C9 5 0 1.00P
R7 5 41 25.0
*
* OUTPUT STAGE
*
Q10 4 41 43 QOUTP1 2.00
Q11 7 41 44 QOUTN1 2.00
Q12 7 43 6 QOUTN2
C15 6 0 1.00P
Q13 4 44 6 QOUTP2
D9 41 6 DY
D10 6 41 DY
*
* NOISE BLOCKS
*
G14 51 50 POLY(1) 14 0 8.09U 4.05U
D11 50 0 DN1
D12 0 51 DN1
*
G15 53 52 POLY(1) 14 0 8.09U 4.05U
D13 52 0 DN2
D14 0 53 DN2
*
G16 55 54 POLY(1) 14 0 2.71U 1.35U
D15 54 0 DN3
D16 0 55 DN3
*
* MODELS
*
.MODEL DN1 D IS=0.166F KF=19.6U AF=3.00
.MODEL DN2 D IS=0.166F KF=18.2U AF=3.00
.MODEL DN3 D IS=0.166F KF=1.07F AF=1.00
.MODEL DX D TT=100N
.MODEL DY D IS=4.11E-16 RS=1.00
.MODEL DZ D IS=3.07E-17 RS=1.00
*
.MODEL QINN1 NPN
+ IS =5.800E-16 BF =3.239E+02  NF =1.000E+00 VAF=4.229E+01
+ IKF=6.700E-02 ISE=8.000E-17  NE =1.197E+00 BR =4.003E+01
+ NR =1.000E+00 VAR=1.696E+00  IKR=1.000E-01 ISC=4.000E-19
+ NC =1.700E+00 RB =1.843E+01  IRB=0.000E+00 RBM=4.083E+00
+ RE =2.100E-01 RC =1.000E+01  CJE=4.300E-13 VJE=7.973E-01
+ MJE=4.950E-01 TF =1.862E-11  XTF=1.873E+01 VTF=2.825E+00
+ ITF=1.651E-01 PTF=0.000E+00  CJC=3.500E-13 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=1.778E-01 TR =7.000E-10 CJS=1.600E-12
+ VJS=5.723E-01 MJS=0.000E+00  FC =9.765E-01
*
.MODEL QINN2 NPN
+ IS =5.800E-16 BF =2.939E+02  NF =1.000E+00 VAF=3.279E+01
+ IKF=6.700E-02 ISE=8.000E-17  NE =1.197E+00 BR =4.003E+01
+ NR =1.000E+00 VAR=1.696E+00  IKR=1.000E-01 ISC=4.000E-19
+ NC =1.700E+00 RB =1.843E+01  IRB=0.000E+00 RBM=4.083E+00
+ RE =2.100E-01 RC =1.000E+01  CJE=4.300E-13 VJE=7.973E-01
+ MJE=4.950E-01 TF =1.862E-11  XTF=1.873E+01 VTF=2.825E+00
+ ITF=1.651E-01 PTF=0.000E+00  CJC=3.500E-13 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=1.778E-01 TR =7.000E-10 CJS=1.600E-12
+ VJS=5.723E-01 MJS=0.000E+00  FC =9.765E-01
*
.MODEL QOUTN1 NPN
+ IS =3.954E-16 BF =3.239E+02  NF =1.000E+00 VAF=8.457E+01
+ IKF=4.590E-02 ISE=5.512E-17  NE =1.197E+00 BR =3.957E+01
+ NR =1.000E+00 VAR=1.696E+00  IKR=7.392E-02 ISC=2.867E-19
+ NC =1.700E+00 RB =3.645E+01  IRB=0.000E+00 RBM=8.077E+00
+ RE =3.010E-01 RC =2.438E+01  CJE=2.962E-13 VJE=7.973E-01
+ MJE=4.950E-01 TF =1.875E-11  XTF=1.873E+01 VTF=2.825E+00
+ ITF=1.110E-01 PTF=0.000E+00  CJC=2.608E-13 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=1.704E-01 TR =5.832E-10 CJS=4.115E-13
+ VJS=5.723E-01 MJS=4.105E-01  FC =9.765E-01
*
.MODEL QOUTN2 NPN
+ IS =1.880E-15 BF =3.239E+02  NF =1.000E+00 VAF=8.457E+01
+ IKF=2.182E-01 ISE=2.620E-16  NE =1.197E+00 BR =4.090E+01
+ NR =1.000E+00 VAR=1.696E+00  IKR=3.513E-01 ISC=1.229E-18
+ NC =1.700E+00 RB =7.668E+00  IRB=0.000E+00 RBM=1.699E+00
+ RE =5.063E+00 RC =3.371E+00  CJE=1.408E-12 VJE=7.973E-01
+ MJE=4.950E-01 TF =1.838E-11  XTF=1.873E+01 VTF=2.825E+00
+ ITF=5.278E-01 PTF=0.000E+00  CJC=1.095E-12 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=1.930E-01 TR =1.296E-09 CJS=1.217E-12
+ VJS=5.723E-01 MJS=4.105E-01  FC =9.765E-01
*
.MODEL QINP1 PNP
+ IS =3.500E-16 BF =7.165E+01  NF =1.000E+00 VAF=1.720E+01
+ IKF=4.120E-02 ISE=1.750E-15  NE =1.366E+00 BR =1.970E+01
+ NR =1.000E+00 VAR=1.805E+00  IKR=3.600E-01 ISC=9.877E-18
+ NC =1.634E+00 RB =7.797E+00  IRB=0.000E+00 RBM=1.915E+00
+ RE =2.260E-01 RC =1.500E+01  CJE=4.300E-13 VJE=7.975E-01
+ MJE=5.000E-01 TF =3.032E-11  XTF=5.386E+00 VTF=2.713E+00
+ ITF=1.374E-01 PTF=0.000E+00  CJC=5.600E-13 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=1.778E-01 TR =1.605E-09 CJS=1.600E-12
+ VJS=6.691E-01 MJS=0.000E+00  FC =8.803E-01
*
.MODEL QINP2 PNP
+ IS =3.500E-16 BF =6.565E+01  NF =1.000E+00 VAF=1.370E+01
+ IKF=4.120E-02 ISE=1.750E-15  NE =1.366E+00 BR =1.970E+01
+ NR =1.000E+00 VAR=1.805E+00  IKR=3.600E-01 ISC=9.877E-18
+ NC =1.634E+00 RB =7.797E+00  IRB=0.000E+00 RBM=1.915E+00
+ RE =2.260E-01 RC =1.500E+01  CJE=4.300E-13 VJE=7.975E-01
+ MJE=5.000E-01 TF =3.032E-11  XTF=5.386E+00 VTF=2.713E+00
+ ITF=1.374E-01 PTF=0.000E+00  CJC=5.600E-13 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=1.778E-01 TR =1.605E-09 CJS=1.600E-12
+ VJS=6.691E-01 MJS=0.000E+00  FC =8.803E-01
*
.MODEL QOUTP1 PNP
+ IS =2.399E-16 BF =7.165E+01  NF =1.000E+00 VAF=3.439E+01
+ IKF=3.509E-02 ISE=1.190E-15  NE =1.366E+00 BR =1.946E+01
+ NR =1.000E+00 VAR=1.805E+00  IKR=2.464E-01 ISC=6.685E-18
+ NC =1.634E+00 RB =1.542E+01  IRB=0.000E+00 RBM=3.788E+00
+ RE =3.281E-01 RC =1.420E+01  CJE=2.962E-13 VJE=7.975E-01
+ MJE=5.000E-01 TF =3.051E-11  XTF=5.386E+00 VTF=2.713E+00
+ ITF=9.481E-02 PTF=0.000E+00  CJC=4.131E-13 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=1.704E-01 TR =1.388E-09 CJS=9.092E-13
+ VJS=6.691E-01 MJS=3.950E-01  FC =8.803E-01
*
.MODEL QOUTP2 PNP
+ IS =1.140E-15 BF =1.401E+02  NF =1.000E+00 VAF=3.439E+01
+ IKF=1.668E-01 ISE=5.655E-15  NE =1.366E+00 BR =2.009E+01
+ NR =1.000E+00 VAR=1.805E+00  IKR=1.171E+00 ISC=3.141E-17
+ NC =1.634E+00 RB =3.245E+00  IRB=0.000E+00 RBM=7.970E-01
+ RE =5.069E+00 RC =5.381E+00  CJE=1.408E-12 VJE=7.975E-01
+ MJE=5.000E-01 TF =3.013E-11  XTF=5.386E+00 VTF=2.713E+00
+ ITF=4.506E-01 PTF=0.000E+00  CJC=1.734E-12 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=1.929E-01 TR =2.704E-09 CJS=2.020E-12
+ VJS=6.691E-01 MJS=3.950E-01  FC =8.803E-01
*
.ENDS 
*$
