
*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Inc.
* Models developed and under copyright by:
* National Semiconductor, Inc.  

*/////////////////////////////////////////////////////////////////////
* Legal Notice: This material is intended for free software support.
* The file may be copied, and distributed; however, reselling the 
*  material is illegal

*////////////////////////////////////////////////////////////////////
* For ordering or technical information on these models, contact:
* National Semiconductor's Customer Response Center
*                 7:00 A.M.--7:00 P.M.  U.S. Central Time
*                                (800) 272-9959
* For Applications support, contact the Internet address:
*  Appshelp@galaxy.nsc.com

*//////////////////////////////////////////////////////////
*LM6310 CURRENT FEEDBACK OP-AMP MACRO-MODEL
*//////////////////////////////////////////////////////////
* Connections:     Non-Inverting Input
*                  | Inverting Input
*                  | | Output
*                  | | | +Vcc
*                  | | | | -Vee
*                  | | | | | Vdis_bar
*                  | | | | | |
.SUBCKT LM6310/NS 3 2 6 7 4 8
*Features
* This is a Low-Cost, Low-Power, 110MHz, Monolithic
* Current Feedback Op Amp with Disable
*
* DISABLE/BIAS BLOCK
*
R1 7 8 20.0K
C3 8 0 1.00P
R2 8 10 5.00K
Q1 7 10 15 QINN
R3 7 12 100
V1 12 13 1.50
Q2 13 14 15 QINN
D1 10 11 DDV
D2 11 10 DDV 0.11
R4 11 14 2.00K
R5 14 16 2.00K
R6 7 16 20.0K
R7 16 17 20.0K
C4 15 0 336F
I1 15 4 150U
C5 17 0 101F
V2 17 4 3.00
*
R8 7 20 20.0K
D3 20 21 DQ 1.88
G1 21 0 POLY(1) 7 12 0 10.0M
D4 22 21 DQ 1.88
Q3 22 20 7 QINP 3.00
I2 22 4 176U
R9 7 23 625
D5 23 22 DDV 0.28
C6 22 0 1.00P
*
C1 7 0 1.00P
C2 4 0 1.00P
G2 7 4 POLY(1) 7 23 0 4.13M
G3 7 30 POLY(1) 7 23 0 1.54M
C7 30 0 751F
G4 34 4 POLY(1) 7 23 0 1.46M
C8 34 0 751F
*
* INPUT STAGE
*
G5 3 0 POLY(3) 7 23 62 0 63 0 0 20.3U 1.00M 1.00M
C9 3 0 1.00P
E1 3 32 POLY(2) 60 0 61 0 -1.50M 1.00 1.00
D6 30 31 DQ 0.25
Q4 4 32 31 QINP
Q5 7 32 33 QINN
D7 33 34 DQ 0.25
G6 41 0 POLY(3) 7 23 64 0 65 0 0 36.4U 1.00M 1.00M
Q6 41 30 42 QINN
D8 42 2 DQ 0.25
C10 2 0 3.50P
D9 2 43 DQ 0.25
Q7 44 34 43 QINP
*
* GAIN STAGE
*
R10 7 40 550
C11 7 40 1.80P
V3 40 41 1.90
C12 41 47 580F
C13 41 51 430F
V4 7 46 750M
D10 51 46 DOR
G7 7 47 POLY(2) 7 40 7 47 0 3.83M 208N
G8 7 51 POLY(1) 7 40 0 9.03M
C14 51 0 950F
*
V5 44 45 1.90
R11 45 4 550
C15 45 4 1.80P
C16 44 47 505F
C17 44 50 270F
D11 48 47 DOR
V6 48 4 1.30
G9 47 4 POLY(2) 45 4 47 4 0 3.91M 2.14U
G10 50 4 POLY(1) 45 4 0 3.18M
C18 50 0 515F
*
* OUTPUT STAGE
*
C19 47 0 904F
Q8 7 47 50 QOUTN1
D12 51 52 DDV 1.67
Q9 4 50 52 QOUTP1
Q10 7 51 6 QOUTN2
C20 6 0 1.00P
C21 6 53 403F
E2 53 0 POLY(2) 3 0 7 23 0 1.00 0 0 -9.09
Q11 4 52 6 QOUTP2
*
* NOISE SOURCES
*
I3 61 60 DC 26.8U
D13 60 0 DN1
D14 0 61 DN1
*
I4 63 62 DC 56.9U
D15 62 0 DN2
D16 0 63 DN2
*
I5 65 64 DC 46.9U
D17 64 0 DN3
D18 0 65 DN3
*
* MODELS
*
.MODEL DDV D IS=0.287F N=2.00 RS=274M CJO=354F M=500M VJ=798M TT=30.4P
.MODEL DN1 D IS=0.166F KF=4.48F AF=1.00
.MODEL DN2 D IS=0.166F KF=20.6F AF=1.00
.MODEL DN3 D IS=0.166F KF=87.6F AF=1.00
.MODEL DOR D TT=100N
.MODEL DQ D IS=0.165F RS=561M CJO=159F M=495M VJ=797M TT=19.2P
*
.MODEL QINN NPN
+ IS =4.242E-17 BF =3.239E+02 NF =1.000E+00 VAF=2.115E+01
+ IKF=6.322E-03 ISE=7.591E-18 NE =1.197E+00 BR =3.355E+01
+ NR =1.000E+00 VAR=1.696E+00 IKR=1.018E-02 ISC=6.091E-20
+ NC =1.700E+00 RB =3.146E+02 IRB=0.000E+00 RBM=1.086E+02
+ RE =2.185E+00 RC =3.022E+01 CJE=4.079E-14 VJE=7.973E-01
+ MJE=4.950E-01 TF =2.078E-11 XTF=1.873E+01 VTF=2.825E+00
+ ITF=1.529E-02 CJC=5.906E-14 VJC=8.046E-01 MJC=4.931E-01
+ XCJC=1.04E-01 TR =1.620E-10 CJS=6.743E-13 MJS=0.000E+00
+ VJS=5.723E-01 FC =9.765E-01
*
.MODEL QOUTN1 NPN
+ IS =2.636E-16 BF =3.239E+02 NF =1.000E+00 VAF=8.457E+01
+ IKF=3.060E-02 ISE=3.674E-17 NE =1.197E+00 BR =3.868E+01
+ NR =1.000E+00 VAR=1.696E+00 IKR=4.928E-02 ISC=2.045E-19
+ NC =1.700E+00 RB =5.467E+01 IRB=0.000E+00 RBM=1.212E+01
+ RE =4.515E-01 RC =1.999E+01 CJE=1.974E-13 VJE=7.973E-01
+ MJE=4.950E-01 TF =1.901E-11 XTF=1.873E+01 VTF=2.825E+00
+ ITF=7.403E-02 CJC=1.883E-13 VJC=8.046E-01 MJC=4.931E-01
+ XCJC=1.57E-01 TR =5.184E-10 CJS=3.540E-13 VJS=5.723E-01
+ MJS=4.105E-01 FC =9.765E-01
*
.MODEL QOUTN2 NPN
+ IS =9.456E-16 BF =3.239E+02 NF =1.000E+00 VAF=8.457E+01
+ IKF=1.098E-01 ISE=1.318E-16 NE =1.197E+00 BR =3.989E+01
+ NR =1.000E+00 VAR=1.696E+00 IKR=1.767E-01 ISC=6.688E-19
+ NC =1.700E+00 RB =6.524E+01 IRB=0.000E+00 RBM=5.338E+01
+ RE =1.013E+01 RC =4.303E+00 CJE=7.082E-13 VJE=7.973E-01
+ MJE=4.950E-01 TF =1.866E-11 XTF=1.873E+01 VTF=2.825E+00
+ ITF=2.655E-01 CJC=6.056E-13 VJC=8.046E-01 MJC=4.931E-01
+ XCJC=1.76E-01 TR =8.748E-10 CJS=8.651E-13 VJS=5.723E-01
+ MJS=4.105E-01 FC =9.765E-01
*
.MODEL QINP PNP
+ IS =4.242E-17 BF =7.165E+01 NF =1.000E+00 VAF=1.720E+01
+ IKF=4.832E-03 ISE=1.639E-16 NE =1.366E+00 BR =1.658E+01
+ NR =1.000E+00 VAR=1.805E+00 IKR=3.394E-02 ISC=9.789E-19
+ NC =1.634E+00 RB =1.620E+02 IRB=0.000E+00 RBM=7.750E+01
+ RE =2.382E+00 RC =3.386E+01 CJE=4.079E-14 VJE=7.975E-01
+ MJE=5.000E-01 TF =3.263E-11 XTF=5.386E+00 VTF=2.713E+00
+ ITF=1.306E-02 CJC=9.356E-14 VJC=7.130E-01 MJC=4.200E-01
+ XCJC=1.04E-01 TR =6.577E-10 CJS=6.743E-13 VJS=6.691E-01
+ MJS=0.000E+00 FC =8.803E-01
*
.MODEL QOUTP1 PNP
+ IS =2.399E-16 BF =7.165E+01 NF =1.000E+00 VAF=3.439E+01
+ IKF=3.509E-02 ISE=1.190E-15 NE =1.366E+00 BR =1.946E+01
+ NR =1.000E+00 VAR=1.805E+00 IKR=2.464E-01 ISC=6.685E-18
+ NC =1.634E+00 RB =1.542E+01 IRB=0.000E+00 RBM=3.788E+00
+ RE =3.281E-01 RC =1.420E+01 CJE=2.962E-13 VJE=7.975E-01
+ MJE=5.000E-01 TF =3.051E-11 XTF=5.386E+00 VTF=2.713E+00
+ ITF=9.481E-02 CJC=4.131E-13 VJC=7.130E-01 MJC=4.200E-01
+ XCJC=1.70E-01 TR =1.388E-09 CJS=9.092E-13 VJS=6.691E-01
+ MJS=3.950E-01 FC =8.803E-01
*
.MODEL QOUTP2 PNP
+ IS =1.147E-15 BF =7.165E+01 NF =1.000E+00 VAF=3.439E+01
+ IKF=1.678E-01 ISE=5.690E-15 NE =1.366E+00 BR =1.961E+01
+ NR =1.000E+00 VAR=1.805E+00 IKR=1.178E+00 ISC=3.188E-17
+ NC =1.634E+00 RB =5.323E+01 IRB=0.000E+00 RBM=5.079E+01
+ RE =1.069E+01 RC =3.177E+00 CJE=1.416E-12 VJE=7.975E-01
+ MJE=5.000E-01 TF =3.042E-11 XTF=5.386E+00 VTF=2.713E+00
+ ITF=4.534E-01 CJC=1.918E-12 VJC=7.130E-01 MJC=4.200E-01
+ XCJC=1.76E-01 TR =1.973E-09 CJS=3.054E-12 VJS=6.691E-01
+ MJS=3.950E-01 FC =8.803E-01
*
.ENDS 
*$
