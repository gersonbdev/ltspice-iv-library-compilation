*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Inc.
* Models developed and under copyright by:
* National Semiconductor, Inc.  

*/////////////////////////////////////////////////////////////////////
* Legal Notice: This material is intended for free software support.
* The file may be copied, and distributed; however, reselling the 
*  material is illegal

*////////////////////////////////////////////////////////////////////
* For ordering or technical information on these models, contact:
* National Semiconductor's Customer Response Center
*                 7:00 A.M.--7:00 P.M.  U.S. Central Time
*                                (800) 272-9959
* For Applications support, contact the Internet address:
*  Appshelp@galaxy.nsc.com

*/////////////////////////////////////////////////
*LM6317 Operational Amplifier Macro-Model
*/////////////////////////////////////////////////
* Connections:     Non-Inverting
*                  |  Inverting
*                  |  |  Output
*                  |  |  |  +Vcc
*                  |  |  |  |  -Vcc
*                  |  |  |  |  |
.SUBCKT LM6317/NS 3  2  6  7  4
*Features
*   This is a High Speed, Unity Gain Stable Monolithic Voltage
*   Feedback Op Amp.

*
* INVERTING BUFFER
*
R1 7 10 318
R2 11 4 214
G1 7 12 POLY(2) 7 4 7 10 -58.71U 19.57U 3.145M
C1 12 0 481F
Q1 11 2 12 QINP
C3 2 0 500F
Q2 10 2 13 QINN
C2 13 0 247F
G2 13 4 POLY(2) 7 4 11 4 -16.66U 5.554U 2.921M
*
R3 7 14 433
V1 14 15 1.62
Q3 15 12 16 QINN
R5 16 21 150
Q4 17 13 16 QINP
V2 17 18 1.57
R4 18 4 433
*
* NON-INVERTING BUFFER
*
R6 7 19 437
V3 19 20 1.64
Q5 20 24 21 QINN
Q6 22 26 21 QINP
V4 22 23 1.62
R7 23 4 437
G3 7 24 POLY(2) 7 4 7 27 -59.29U 19.43U 3.145M
C5 24 0 481F
Q7 28 25 24 QINP
C4 25 0 500F
Q8 27 25 26 QINN
C6 26 0 247F
G4 26 4 POLY(2) 7 4 28 4 -17.09U 5.697U 2.912M
R8 7 27 318
E1 3 25 POLY(1) 40 0 500U 2.49
G5 3 0 POLY(1) 41 0 180N 262U
R9 28 4 214
*
* CURRENT MIRROR GAIN BLOCKS
*
V5 7 29 2.10
D1 31 29 DX
C7 20 31 431F
C8 20 6 1.80P
C9 22 6 1.80P
C10 22 31 476F
D2 30 31 DX
V6 30 4 2.10
G6 7 31 POLY(1) 7 19 0 6.865M
R10 31 0 167K
C11 31 0 475F
G7 31 4 POLY(1) 23 4 0 6.865M
G8 7 32 POLY(1) 7 19 0 2.288M
C12 32 0 1.5P
G9 35 4 POLY(1) 23 4 0 2.288M
C13 35 0 1.5P
*
* OUTPUT STAGE
*
D3 32 33 DY
Q9 4 31 33 QOUTP1
Q10 7 31 34 QOUTN1
D4 34 35 DY
Q11 7 32 36 QOUTN1
Q12 4 31 36 QOUTP1
Q13 7 31 37 QOUTN1
Q14 4 35 37 QOUTP1
Q15 7 36 38 QOUTN2
R11 38 6 10.0
C14 6 0 3.20P
R12 6 39 10.0
Q16 4 37 39 QOUTP2
*
* NOISE BLOCKS
*
R13 40 0 122
R14 40 0 122
R15 41 0 122
R16 41 0 122
*
* MODELS
*
.Model DX D TT=200N
.Model DY D IS=0.395F
.Model DZ D IS=0.240F
*
.MODEL QINN NPN
+ IS =0.166F    BF =3.239E+02 NF =1.000E+00 VAF=8.457E+01
+ IKF=2.462E-02 ISE=2.956E-17 NE =1.197E+00 BR =3.719E+01
+ NR =1.000E+00 VAR=1.696E+00 IKR=3.964E-02 ISC=1.835E-19
+ NC =1.700E+00 RB =118       IRB=0.000E+00 RBM=65.1
+ RC =2.645E+01 CJE=1.632E-13 VJE=7.973E-01
+ MJE=4.950E-01 TF =1.948E-11 XTF=1.873E+01 VTF=2.825E+00
+ ITF=5.955E-02 PTF=0.000E+00 CJC=1.720E-13 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=589M     TR =4.212E-10 CJS=629F
+ MJS=0         KF =1.00P     AF =1.000E+00
+ FC =9.765E-01
*
.MODEL QOUTN1 NPN
+ IS =3.954E-16 BF =3.239E+02  NF =1.000E+00 VAF=8.457E+01
+ IKF=4.590E-02 ISE=5.512E-17  NE =1.197E+00 BR =3.719E+01
+ NR =1.000E+00 VAR=1.696E+00  IKR=7.392E-02 ISC=3.087E-19
+ NC =1.700E+00 RB =3.645E+01  IRB=0.000E+00 RBM=8.077E+00
+ RC =2.702E+01 CJE=2.962E-13  VJE=7.973E-01
+ MJE=4.950E-01 TF =1.904E-11  XTF=1.873E+01 VTF=2.825E+00
+ ITF=1.110E-01 PTF=0.000E+00  CJC=2.846E-13 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=1.562E-01 TR =5.832E-10 CJS=5.015E-13
+ VJS=5.723E-01 MJS=4.105E-01  KF =1.00P     AF =1.000E+00
+ FC =9.765E-01
*
.MODEL QOUTN2 NPN
+ IS =9.386E-16 BF =3.239E+02 NF =1.000E+00 VAF=8.457E+01
+ IKF=1.089E-01 ISE=1.308E-16 NE =1.197E+00 BR =3.960E+01
+ NR =1.000E+00 VAR=1.696E+00 IKR=1.754E-01 ISC=6.787E-19
+ NC =1.700E+00 RB =15.4      IRB=0.000E+00 RBM=3.4
+ RC =1.857E+01 CJE=7.030E-13 VJE=7.973E-01
+ MJE=4.950E-01 TF =1.874E-11 XTF=1.873E+01 VTF=2.825E+00
+ ITF=2.635E-01 PTF=0.000E+00 CJC=6.172E-13 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=171M     TR =1.069E-09 CJS=1.028E-12
+ VJS=5.723E-01 MJS=4.105E-01 KF =1.00P     AF =1.000E+00
+ FC =9.765E-01
*
.MODEL QINP PNP
+ IS =0.166F    BF =7.165E+01 NF =1.000E+00 VAF=20.0
+ IKF=1.882E-02 ISE=6.380E-16 NE =1.366E+00 BR =1.833E+01
+ NR =1.000E+00 VAR=1.805E+00 IKR=1.321E-01 ISC=3.666E-18
+ NC =1.634E+00 RB =78.8      IRB=0.000E+00 RBM=57.6
+ RC =3.739E+01 CJE=1.588E-13 VJE=7.975E-01
+ MJE=5.000E-01 TF =3.156E-11 XTF=5.386E+00 VTF=2.713E+00
+ ITF=5.084E-02 PTF=0.000E+00 CJC=2.725E-13 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=741M     TR =7.500E-11 CJS=515F
+ MJS=0         KF =1.00P     AF =1.000E+00
+ FC =8.803E-01
*
.MODEL QOUTP1 PNP
+ IS =2.399E-16 BF =7.165E+01  NF =1.000E+00 VAF=3.439E+01
+ IKF=3.509E-02 ISE=1.190E-15  NE =1.366E+00 BR =1.900E+01
+ NR =1.000E+00 VAR=1.805E+00  IKR=2.464E-01 ISC=6.745E-18
+ NC =1.634E+00 RB =1.542E+01  IRB=0.000E+00 RBM=4.059E+00
+ RC =4.174E+01 CJE=2.962E-13  VJE=7.975E-01
+ MJE=5.000E-01 TF =3.107E-11  XTF=5.386E+00 VTF=2.713E+00
+ ITF=9.481E-02 PTF=0.000E+00  CJC=4.508E-13 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=1.562E-01 TR =9.500E-11 CJS=1.045E-12
+ VJS=6.691E-01 MJS=3.950E-01  KF =1.00P     AF =1.000E+00
+ FC =8.803E-01
*
.MODEL QOUTP2 PNP
+ IS =5.693E-16 BF =7.165E+01 NF =1.000E+00 VAF=3.439E+01
+ IKF=8.328E-02 ISE=2.824E-15 NE =1.366E+00 BR =1.948E+01
+ NR =1.000E+00 VAR=1.805E+00 IKR=5.848E-01 ISC=1.586E-17
+ NC =1.634E+00 RB =6.5       IRB=0.000E+00 RBM=1.7
+ RC =1.767E+01 CJE=7.030E-13 VJE=7.975E-01
+ MJE=5.000E-01 TF =3.073E-11 XTF=5.386E+00 VTF=2.713E+00
+ ITF=2.250E-01 PTF=0.000E+00 CJC=9.776E-13 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=171M     TR =1.450E-10 CJS=1.637E-12
+ VJS=6.691E-01 MJS=3.950E-01 KF =1.00P     AF =1.000E+00
+ FC =8.803E-01
*
.ENDS
 *$
